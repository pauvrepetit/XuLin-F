   
    parameter PROC_NUM = 35;
    parameter ST_IDLE = 3'b000;
    parameter ST_FILTER_FAKE = 3'b001;
    parameter ST_DL_DETECTED = 3'b010;
    parameter ST_DL_REPORT = 3'b100;
   

    reg [2:0] CS_fsm;
    reg [2:0] NS_fsm;
    reg [PROC_NUM - 1:0] dl_detect_reg;
    reg [PROC_NUM - 1:0] dl_done_reg;
    reg [PROC_NUM - 1:0] origin_reg;
    reg [PROC_NUM - 1:0] dl_in_vec_reg;
    reg [31:0] dl_keep_cnt;
    integer i;
    integer fp;

    // FSM State machine
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            CS_fsm <= ST_IDLE;
        end
        else begin
            CS_fsm <= NS_fsm;
        end
    end
    always @ (CS_fsm or dl_in_vec or dl_detect_reg or dl_done_reg or dl_in_vec or origin_reg or dl_keep_cnt) begin
        case (CS_fsm)
            ST_IDLE : begin
                if (|dl_in_vec) begin
                    NS_fsm = ST_FILTER_FAKE;
                end
                else begin
                    NS_fsm = ST_IDLE;
                end
            end
            ST_FILTER_FAKE: begin
                if (dl_keep_cnt >= 32'd1000) begin
                    NS_fsm = ST_DL_DETECTED;
                end
                else if (dl_detect_reg != (dl_detect_reg & dl_in_vec)) begin
                    NS_fsm = ST_IDLE;
                end
                else begin
                    NS_fsm = ST_FILTER_FAKE;
                end
            end
            ST_DL_DETECTED: begin
                // has unreported deadlock cycle
                if (dl_detect_reg != dl_done_reg) begin
                    NS_fsm = ST_DL_REPORT;
                end
                else begin
                    NS_fsm = ST_DL_DETECTED;
                end
            end
            ST_DL_REPORT: begin
                if (|(dl_in_vec & origin_reg)) begin
                    NS_fsm = ST_DL_DETECTED;
                end
                else begin
                    NS_fsm = ST_DL_REPORT;
                end
            end
            default: NS_fsm = ST_IDLE;
        endcase
    end

    // dl_detect_reg record the procs that first detect deadlock
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            dl_detect_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_IDLE) begin
                dl_detect_reg <= dl_in_vec;
            end
        end
    end

    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            dl_keep_cnt <= 32'h0;
        end
        else begin
            if (CS_fsm == ST_FILTER_FAKE && (dl_detect_reg == (dl_detect_reg & dl_in_vec))) begin
                dl_keep_cnt <= dl_keep_cnt + 32'h1;
            end
            else if (CS_fsm == ST_FILTER_FAKE && (dl_detect_reg != (dl_detect_reg & dl_in_vec))) begin
                dl_keep_cnt <= 32'h0;
            end
        end
    end

    // dl_detect_out keeps in high after deadlock detected
    assign dl_detect_out = (|dl_detect_reg) && (CS_fsm == ST_DL_DETECTED || CS_fsm == ST_DL_REPORT);

    // dl_done_reg record the cycles has been reported
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            dl_done_reg <= 'b0;
        end
        else begin
            if ((CS_fsm == ST_DL_REPORT) && (|(dl_in_vec & dl_detect_reg) == 'b1)) begin
                dl_done_reg <= dl_done_reg | dl_in_vec;
            end
        end
    end

    // clear token once a cycle is done
    assign token_clear = (CS_fsm == ST_DL_REPORT) ? ((|(dl_in_vec & origin_reg)) ? 'b1 : 'b0) : 'b0;

    // origin_reg record the current cycle start id
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            origin_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED) begin
                origin_reg <= origin;
            end
        end
    end
   
    // origin will be valid for only one cycle
    wire [PROC_NUM*PROC_NUM - 1:0] origin_tmp;
    assign origin_tmp[PROC_NUM - 1:0] = (dl_detect_reg[0] & ~dl_done_reg[0]) ? 'b1 : 'b0;
    genvar j;
    generate
    for(j = 1;j < PROC_NUM;j = j + 1) begin: F1
        assign origin_tmp[j*PROC_NUM +: PROC_NUM] = (dl_detect_reg[j] & ~dl_done_reg[j]) ? ('b1 << j) : origin_tmp[(j - 1)*PROC_NUM +: PROC_NUM];
    end
    endgenerate
    always @ (CS_fsm or origin_tmp) begin
        if (CS_fsm == ST_DL_DETECTED) begin
            origin = origin_tmp[(PROC_NUM - 1)*PROC_NUM +: PROC_NUM];
        end
        else begin
            origin = 'b0;
        end
    end

    
    // dl_in_vec_reg record the current cycle dl_in_vec
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            dl_in_vec_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED) begin
                dl_in_vec_reg <= origin;
            end
            else if (CS_fsm == ST_DL_REPORT) begin
                dl_in_vec_reg <= dl_in_vec;
            end
        end
    end
    
    // find_df_deadlock to report the deadlock
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            find_df_deadlock <= 1'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED && dl_detect_reg == dl_done_reg) begin
                find_df_deadlock <= 1'b1;
            end
            else if (CS_fsm == ST_IDLE) begin
                find_df_deadlock <= 1'b0;
            end
        end
    end
    
    // get the first valid proc index in dl vector
    function integer proc_index(input [PROC_NUM - 1:0] dl_vec);
        begin
            proc_index = 0;
            for (i = 0; i < PROC_NUM; i = i + 1) begin
                if (dl_vec[i]) begin
                    proc_index = i;
                end
            end
        end
    endfunction

    // get the proc path based on dl vector
    function [336:0] proc_path(input [PROC_NUM - 1:0] dl_vec);
        integer index;
        begin
            index = proc_index(dl_vec);
            case (index)
                0 : begin
                    proc_path = "kernel_pr_kernel_pr.entry_proc_U0";
                end
                1 : begin
                    proc_path = "kernel_pr_kernel_pr.load_bipedge_U0";
                end
                2 : begin
                    proc_path = "kernel_pr_kernel_pr.load_bipedge_1_U0";
                end
                3 : begin
                    proc_path = "kernel_pr_kernel_pr.load_value_U0";
                end
                4 : begin
                    proc_path = "kernel_pr_kernel_pr.load_value_1_U0";
                end
                5 : begin
                    proc_path = "kernel_pr_kernel_pr.load_value_2_U0";
                end
                6 : begin
                    proc_path = "kernel_pr_kernel_pr.load_value_3_U0";
                end
                7 : begin
                    proc_path = "kernel_pr_kernel_pr.load_value_4_U0";
                end
                8 : begin
                    proc_path = "kernel_pr_kernel_pr.load_value_5_U0";
                end
                9 : begin
                    proc_path = "kernel_pr_kernel_pr.load_value_6_U0";
                end
                10 : begin
                    proc_path = "kernel_pr_kernel_pr.load_value_7_U0";
                end
                11 : begin
                    proc_path = "kernel_pr_kernel_pr.load_value_8_U0";
                end
                12 : begin
                    proc_path = "kernel_pr_kernel_pr.load_value_9_U0";
                end
                13 : begin
                    proc_path = "kernel_pr_kernel_pr.load_value_10_U0";
                end
                14 : begin
                    proc_path = "kernel_pr_kernel_pr.load_value_11_U0";
                end
                15 : begin
                    proc_path = "kernel_pr_kernel_pr.load_value_12_U0";
                end
                16 : begin
                    proc_path = "kernel_pr_kernel_pr.load_value_13_U0";
                end
                17 : begin
                    proc_path = "kernel_pr_kernel_pr.load_value_14_U0";
                end
                18 : begin
                    proc_path = "kernel_pr_kernel_pr.load_value_15_U0";
                end
                19 : begin
                    proc_path = "kernel_pr_kernel_pr.write_back_U0";
                end
                20 : begin
                    proc_path = "kernel_pr_kernel_pr.write_back_1_U0";
                end
                21 : begin
                    proc_path = "kernel_pr_kernel_pr.write_back_2_U0";
                end
                22 : begin
                    proc_path = "kernel_pr_kernel_pr.write_back_3_U0";
                end
                23 : begin
                    proc_path = "kernel_pr_kernel_pr.write_back_4_U0";
                end
                24 : begin
                    proc_path = "kernel_pr_kernel_pr.write_back_5_U0";
                end
                25 : begin
                    proc_path = "kernel_pr_kernel_pr.write_back_6_U0";
                end
                26 : begin
                    proc_path = "kernel_pr_kernel_pr.write_back_7_U0";
                end
                27 : begin
                    proc_path = "kernel_pr_kernel_pr.write_back_8_U0";
                end
                28 : begin
                    proc_path = "kernel_pr_kernel_pr.write_back_9_U0";
                end
                29 : begin
                    proc_path = "kernel_pr_kernel_pr.write_back_10_U0";
                end
                30 : begin
                    proc_path = "kernel_pr_kernel_pr.write_back_11_U0";
                end
                31 : begin
                    proc_path = "kernel_pr_kernel_pr.write_back_12_U0";
                end
                32 : begin
                    proc_path = "kernel_pr_kernel_pr.write_back_13_U0";
                end
                33 : begin
                    proc_path = "kernel_pr_kernel_pr.write_back_14_U0";
                end
                34 : begin
                    proc_path = "kernel_pr_kernel_pr.write_back_15_U0";
                end
                default : begin
                    proc_path = "unknown";
                end
            endcase
        end
    endfunction

    // print the headlines of deadlock detection
    task print_dl_head;
        begin
            $display("\n//////////////////////////////////////////////////////////////////////////////");
            $display("// ERROR!!! DEADLOCK DETECTED at %0t ns! SIMULATION WILL BE STOPPED! //", $time);
            $display("//////////////////////////////////////////////////////////////////////////////");
            fp = $fopen("deadlock_db.dat", "w");
        end
    endtask

    // print the start of a cycle
    task print_cycle_start(input reg [336:0] proc_path, input integer cycle_id);
        begin
            $display("/////////////////////////");
            $display("// Dependence cycle %0d:", cycle_id);
            $display("// (1): Process: %0s", proc_path);
            $fdisplay(fp, "Dependence_Cycle_ID %0d", cycle_id);
            $fdisplay(fp, "Dependence_Process_ID 1");
            $fdisplay(fp, "Dependence_Process_path %0s", proc_path);
        end
    endtask

    // print the end of deadlock detection
    task print_dl_end(input integer num, input integer record_time);
        begin
            $display("////////////////////////////////////////////////////////////////////////");
            $display("// Totally %0d cycles detected!", num);
            $display("////////////////////////////////////////////////////////////////////////");
            $display("// ERROR!!! DEADLOCK DETECTED at %0t ns! SIMULATION WILL BE STOPPED! //", record_time);
            $display("//////////////////////////////////////////////////////////////////////////////");
            $fdisplay(fp, "Dependence_Cycle_Number %0d", num);
            $fclose(fp);
        end
    endtask

    // print one proc component in the cycle
    task print_cycle_proc_comp(input reg [336:0] proc_path, input integer cycle_comp_id);
        begin
            $display("// (%0d): Process: %0s", cycle_comp_id, proc_path);
            $fdisplay(fp, "Dependence_Process_ID %0d", cycle_comp_id);
            $fdisplay(fp, "Dependence_Process_path %0s", proc_path);
        end
    endtask

    // print one channel component in the cycle
    task print_cycle_chan_comp(input [PROC_NUM - 1:0] dl_vec1, input [PROC_NUM - 1:0] dl_vec2);
        reg [424:0] chan_path;
        integer index1;
        integer index2;
        begin
            index1 = proc_index(dl_vec1);
            index2 = proc_index(dl_vec2);
            case (index1)
                0 : begin
                    case(index2)
                    19: begin
                        if (~entry_proc_U0.H_write0_c_blk_n) begin
                            if (~H_write0_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write0_c_U' written by process 'kernel_pr_kernel_pr.write_back_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write0_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write0_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write0_c_U' read by process 'kernel_pr_kernel_pr.write_back_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write0_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~entry_proc_U0.hyperedge_size_c85_blk_n) begin
                            if (~hyperedge_size_c85_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c85_U' written by process 'kernel_pr_kernel_pr.write_back_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c85_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c85_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c85_U' read by process 'kernel_pr_kernel_pr.write_back_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c85_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back_U0_U.if_full_n & entry_proc_U0.ap_start & ~entry_proc_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back_U0_U' read by process 'kernel_pr_kernel_pr.write_back_U0',");
                        end
                    end
                    20: begin
                        if (~entry_proc_U0.H_write1_c_blk_n) begin
                            if (~H_write1_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write1_c_U' written by process 'kernel_pr_kernel_pr.write_back_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write1_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write1_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write1_c_U' read by process 'kernel_pr_kernel_pr.write_back_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write1_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~entry_proc_U0.hyperedge_size_c84_blk_n) begin
                            if (~hyperedge_size_c84_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c84_U' written by process 'kernel_pr_kernel_pr.write_back_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c84_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c84_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c84_U' read by process 'kernel_pr_kernel_pr.write_back_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c84_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back_1_U0_U.if_full_n & entry_proc_U0.ap_start & ~entry_proc_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back_1_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back_1_U0_U' read by process 'kernel_pr_kernel_pr.write_back_1_U0',");
                        end
                    end
                    21: begin
                        if (~entry_proc_U0.H_write2_c_blk_n) begin
                            if (~H_write2_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write2_c_U' written by process 'kernel_pr_kernel_pr.write_back_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write2_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write2_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write2_c_U' read by process 'kernel_pr_kernel_pr.write_back_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write2_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~entry_proc_U0.hyperedge_size_c83_blk_n) begin
                            if (~hyperedge_size_c83_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c83_U' written by process 'kernel_pr_kernel_pr.write_back_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c83_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c83_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c83_U' read by process 'kernel_pr_kernel_pr.write_back_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c83_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back_2_U0_U.if_full_n & entry_proc_U0.ap_start & ~entry_proc_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back_2_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back_2_U0_U' read by process 'kernel_pr_kernel_pr.write_back_2_U0',");
                        end
                    end
                    22: begin
                        if (~entry_proc_U0.H_write3_c_blk_n) begin
                            if (~H_write3_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write3_c_U' written by process 'kernel_pr_kernel_pr.write_back_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write3_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write3_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write3_c_U' read by process 'kernel_pr_kernel_pr.write_back_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write3_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~entry_proc_U0.hyperedge_size_c82_blk_n) begin
                            if (~hyperedge_size_c82_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c82_U' written by process 'kernel_pr_kernel_pr.write_back_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c82_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c82_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c82_U' read by process 'kernel_pr_kernel_pr.write_back_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c82_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back_3_U0_U.if_full_n & entry_proc_U0.ap_start & ~entry_proc_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back_3_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back_3_U0_U' read by process 'kernel_pr_kernel_pr.write_back_3_U0',");
                        end
                    end
                    23: begin
                        if (~entry_proc_U0.H_write4_c_blk_n) begin
                            if (~H_write4_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write4_c_U' written by process 'kernel_pr_kernel_pr.write_back_4_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write4_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write4_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write4_c_U' read by process 'kernel_pr_kernel_pr.write_back_4_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write4_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~entry_proc_U0.hyperedge_size_c81_blk_n) begin
                            if (~hyperedge_size_c81_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c81_U' written by process 'kernel_pr_kernel_pr.write_back_4_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c81_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c81_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c81_U' read by process 'kernel_pr_kernel_pr.write_back_4_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c81_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back_4_U0_U.if_full_n & entry_proc_U0.ap_start & ~entry_proc_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back_4_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back_4_U0_U' read by process 'kernel_pr_kernel_pr.write_back_4_U0',");
                        end
                    end
                    24: begin
                        if (~entry_proc_U0.H_write5_c_blk_n) begin
                            if (~H_write5_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write5_c_U' written by process 'kernel_pr_kernel_pr.write_back_5_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write5_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write5_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write5_c_U' read by process 'kernel_pr_kernel_pr.write_back_5_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write5_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~entry_proc_U0.hyperedge_size_c80_blk_n) begin
                            if (~hyperedge_size_c80_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c80_U' written by process 'kernel_pr_kernel_pr.write_back_5_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c80_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c80_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c80_U' read by process 'kernel_pr_kernel_pr.write_back_5_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c80_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back_5_U0_U.if_full_n & entry_proc_U0.ap_start & ~entry_proc_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back_5_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back_5_U0_U' read by process 'kernel_pr_kernel_pr.write_back_5_U0',");
                        end
                    end
                    25: begin
                        if (~entry_proc_U0.H_write6_c_blk_n) begin
                            if (~H_write6_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write6_c_U' written by process 'kernel_pr_kernel_pr.write_back_6_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write6_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write6_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write6_c_U' read by process 'kernel_pr_kernel_pr.write_back_6_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write6_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~entry_proc_U0.hyperedge_size_c79_blk_n) begin
                            if (~hyperedge_size_c79_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c79_U' written by process 'kernel_pr_kernel_pr.write_back_6_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c79_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c79_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c79_U' read by process 'kernel_pr_kernel_pr.write_back_6_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c79_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back_6_U0_U.if_full_n & entry_proc_U0.ap_start & ~entry_proc_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back_6_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back_6_U0_U' read by process 'kernel_pr_kernel_pr.write_back_6_U0',");
                        end
                    end
                    26: begin
                        if (~entry_proc_U0.H_write7_c_blk_n) begin
                            if (~H_write7_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write7_c_U' written by process 'kernel_pr_kernel_pr.write_back_7_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write7_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write7_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write7_c_U' read by process 'kernel_pr_kernel_pr.write_back_7_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write7_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~entry_proc_U0.hyperedge_size_c78_blk_n) begin
                            if (~hyperedge_size_c78_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c78_U' written by process 'kernel_pr_kernel_pr.write_back_7_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c78_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c78_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c78_U' read by process 'kernel_pr_kernel_pr.write_back_7_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c78_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back_7_U0_U.if_full_n & entry_proc_U0.ap_start & ~entry_proc_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back_7_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back_7_U0_U' read by process 'kernel_pr_kernel_pr.write_back_7_U0',");
                        end
                    end
                    27: begin
                        if (~entry_proc_U0.H_write8_c_blk_n) begin
                            if (~H_write8_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write8_c_U' written by process 'kernel_pr_kernel_pr.write_back_8_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write8_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write8_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write8_c_U' read by process 'kernel_pr_kernel_pr.write_back_8_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write8_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~entry_proc_U0.hyperedge_size_c77_blk_n) begin
                            if (~hyperedge_size_c77_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c77_U' written by process 'kernel_pr_kernel_pr.write_back_8_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c77_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c77_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c77_U' read by process 'kernel_pr_kernel_pr.write_back_8_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c77_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back_8_U0_U.if_full_n & entry_proc_U0.ap_start & ~entry_proc_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back_8_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back_8_U0_U' read by process 'kernel_pr_kernel_pr.write_back_8_U0',");
                        end
                    end
                    28: begin
                        if (~entry_proc_U0.H_write9_c_blk_n) begin
                            if (~H_write9_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write9_c_U' written by process 'kernel_pr_kernel_pr.write_back_9_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write9_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write9_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write9_c_U' read by process 'kernel_pr_kernel_pr.write_back_9_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write9_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~entry_proc_U0.hyperedge_size_c76_blk_n) begin
                            if (~hyperedge_size_c76_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c76_U' written by process 'kernel_pr_kernel_pr.write_back_9_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c76_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c76_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c76_U' read by process 'kernel_pr_kernel_pr.write_back_9_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c76_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back_9_U0_U.if_full_n & entry_proc_U0.ap_start & ~entry_proc_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back_9_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back_9_U0_U' read by process 'kernel_pr_kernel_pr.write_back_9_U0',");
                        end
                    end
                    29: begin
                        if (~entry_proc_U0.H_write10_c_blk_n) begin
                            if (~H_write10_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write10_c_U' written by process 'kernel_pr_kernel_pr.write_back_10_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write10_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write10_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write10_c_U' read by process 'kernel_pr_kernel_pr.write_back_10_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write10_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~entry_proc_U0.hyperedge_size_c75_blk_n) begin
                            if (~hyperedge_size_c75_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c75_U' written by process 'kernel_pr_kernel_pr.write_back_10_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c75_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c75_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c75_U' read by process 'kernel_pr_kernel_pr.write_back_10_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c75_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back_10_U0_U.if_full_n & entry_proc_U0.ap_start & ~entry_proc_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back_10_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back_10_U0_U' read by process 'kernel_pr_kernel_pr.write_back_10_U0',");
                        end
                    end
                    30: begin
                        if (~entry_proc_U0.H_write11_c_blk_n) begin
                            if (~H_write11_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write11_c_U' written by process 'kernel_pr_kernel_pr.write_back_11_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write11_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write11_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write11_c_U' read by process 'kernel_pr_kernel_pr.write_back_11_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write11_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~entry_proc_U0.hyperedge_size_c74_blk_n) begin
                            if (~hyperedge_size_c74_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c74_U' written by process 'kernel_pr_kernel_pr.write_back_11_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c74_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c74_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c74_U' read by process 'kernel_pr_kernel_pr.write_back_11_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c74_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back_11_U0_U.if_full_n & entry_proc_U0.ap_start & ~entry_proc_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back_11_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back_11_U0_U' read by process 'kernel_pr_kernel_pr.write_back_11_U0',");
                        end
                    end
                    31: begin
                        if (~entry_proc_U0.H_write12_c_blk_n) begin
                            if (~H_write12_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write12_c_U' written by process 'kernel_pr_kernel_pr.write_back_12_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write12_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write12_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write12_c_U' read by process 'kernel_pr_kernel_pr.write_back_12_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write12_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~entry_proc_U0.hyperedge_size_c73_blk_n) begin
                            if (~hyperedge_size_c73_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c73_U' written by process 'kernel_pr_kernel_pr.write_back_12_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c73_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c73_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c73_U' read by process 'kernel_pr_kernel_pr.write_back_12_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c73_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back_12_U0_U.if_full_n & entry_proc_U0.ap_start & ~entry_proc_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back_12_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back_12_U0_U' read by process 'kernel_pr_kernel_pr.write_back_12_U0',");
                        end
                    end
                    32: begin
                        if (~entry_proc_U0.H_write13_c_blk_n) begin
                            if (~H_write13_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write13_c_U' written by process 'kernel_pr_kernel_pr.write_back_13_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write13_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write13_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write13_c_U' read by process 'kernel_pr_kernel_pr.write_back_13_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write13_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~entry_proc_U0.hyperedge_size_c72_blk_n) begin
                            if (~hyperedge_size_c72_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c72_U' written by process 'kernel_pr_kernel_pr.write_back_13_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c72_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c72_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c72_U' read by process 'kernel_pr_kernel_pr.write_back_13_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c72_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back_13_U0_U.if_full_n & entry_proc_U0.ap_start & ~entry_proc_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back_13_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back_13_U0_U' read by process 'kernel_pr_kernel_pr.write_back_13_U0',");
                        end
                    end
                    33: begin
                        if (~entry_proc_U0.H_write14_c_blk_n) begin
                            if (~H_write14_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write14_c_U' written by process 'kernel_pr_kernel_pr.write_back_14_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write14_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write14_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write14_c_U' read by process 'kernel_pr_kernel_pr.write_back_14_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write14_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~entry_proc_U0.hyperedge_size_c71_blk_n) begin
                            if (~hyperedge_size_c71_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c71_U' written by process 'kernel_pr_kernel_pr.write_back_14_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c71_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c71_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c71_U' read by process 'kernel_pr_kernel_pr.write_back_14_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c71_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back_14_U0_U.if_full_n & entry_proc_U0.ap_start & ~entry_proc_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back_14_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back_14_U0_U' read by process 'kernel_pr_kernel_pr.write_back_14_U0',");
                        end
                    end
                    34: begin
                        if (~entry_proc_U0.H_write15_c_blk_n) begin
                            if (~H_write15_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write15_c_U' written by process 'kernel_pr_kernel_pr.write_back_15_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write15_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write15_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write15_c_U' read by process 'kernel_pr_kernel_pr.write_back_15_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write15_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~entry_proc_U0.hyperedge_size_c_blk_n) begin
                            if (~hyperedge_size_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c_U' written by process 'kernel_pr_kernel_pr.write_back_15_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c_U' read by process 'kernel_pr_kernel_pr.write_back_15_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back_15_U0_U.if_full_n & entry_proc_U0.ap_start & ~entry_proc_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back_15_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back_15_U0_U' read by process 'kernel_pr_kernel_pr.write_back_15_U0',");
                        end
                    end
                    1: begin
                        if (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_load_bipedge_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge_U0'");
                        end
                    end
                    2: begin
                        if (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_load_bipedge_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge_1_U0'");
                        end
                    end
                    3: begin
                        if (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_load_value_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_U0'");
                        end
                    end
                    4: begin
                        if (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_load_value_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_1_U0'");
                        end
                    end
                    5: begin
                        if (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_load_value_2_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_2_U0'");
                        end
                    end
                    6: begin
                        if (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_load_value_3_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_3_U0'");
                        end
                    end
                    7: begin
                        if (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_load_value_4_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_4_U0'");
                        end
                    end
                    8: begin
                        if (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_load_value_5_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_5_U0'");
                        end
                    end
                    9: begin
                        if (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_load_value_6_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_6_U0'");
                        end
                    end
                    10: begin
                        if (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_load_value_7_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_7_U0'");
                        end
                    end
                    11: begin
                        if (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_load_value_8_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_8_U0'");
                        end
                    end
                    12: begin
                        if (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_load_value_9_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_9_U0'");
                        end
                    end
                    13: begin
                        if (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_load_value_10_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_10_U0'");
                        end
                    end
                    14: begin
                        if (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_load_value_11_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_11_U0'");
                        end
                    end
                    15: begin
                        if (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_load_value_12_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_12_U0'");
                        end
                    end
                    16: begin
                        if (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_load_value_13_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_13_U0'");
                        end
                    end
                    17: begin
                        if (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_load_value_14_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_14_U0'");
                        end
                    end
                    18: begin
                        if (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_load_value_15_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_15_U0'");
                        end
                    end
                    endcase
                end
                1 : begin
                    case(index2)
                    3: begin
                        if (~load_bipedge_U0.grp_load_bipedge_Pipeline_load_bipedge_loop_fu_86.bipedge_stream_0_blk_n) begin
                            if (~bipedge_stream_0_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_0_U' written by process 'kernel_pr_kernel_pr.load_value_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_0_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_0_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_0_U' read by process 'kernel_pr_kernel_pr.load_value_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_0_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_bipedge_U0_ap_ready & load_bipedge_U0.ap_idle & ~ap_sync_load_value_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_U0'");
                        end
                    end
                    4: begin
                        if (~load_bipedge_U0.grp_load_bipedge_Pipeline_load_bipedge_loop_fu_86.bipedge_stream_1_blk_n) begin
                            if (~bipedge_stream_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_1_U' written by process 'kernel_pr_kernel_pr.load_value_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_1_U' read by process 'kernel_pr_kernel_pr.load_value_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_bipedge_U0_ap_ready & load_bipedge_U0.ap_idle & ~ap_sync_load_value_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_1_U0'");
                        end
                    end
                    5: begin
                        if (~load_bipedge_U0.grp_load_bipedge_Pipeline_load_bipedge_loop_fu_86.bipedge_stream_2_blk_n) begin
                            if (~bipedge_stream_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_2_U' written by process 'kernel_pr_kernel_pr.load_value_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_2_U' read by process 'kernel_pr_kernel_pr.load_value_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_bipedge_U0_ap_ready & load_bipedge_U0.ap_idle & ~ap_sync_load_value_2_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_2_U0'");
                        end
                    end
                    6: begin
                        if (~load_bipedge_U0.grp_load_bipedge_Pipeline_load_bipedge_loop_fu_86.bipedge_stream_3_blk_n) begin
                            if (~bipedge_stream_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_3_U' written by process 'kernel_pr_kernel_pr.load_value_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_3_U' read by process 'kernel_pr_kernel_pr.load_value_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_bipedge_U0_ap_ready & load_bipedge_U0.ap_idle & ~ap_sync_load_value_3_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_3_U0'");
                        end
                    end
                    7: begin
                        if (~load_bipedge_U0.grp_load_bipedge_Pipeline_load_bipedge_loop_fu_86.bipedge_stream_4_blk_n) begin
                            if (~bipedge_stream_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_4_U' written by process 'kernel_pr_kernel_pr.load_value_4_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_4_U' read by process 'kernel_pr_kernel_pr.load_value_4_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_bipedge_U0_ap_ready & load_bipedge_U0.ap_idle & ~ap_sync_load_value_4_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_4_U0'");
                        end
                    end
                    8: begin
                        if (~load_bipedge_U0.grp_load_bipedge_Pipeline_load_bipedge_loop_fu_86.bipedge_stream_5_blk_n) begin
                            if (~bipedge_stream_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_5_U' written by process 'kernel_pr_kernel_pr.load_value_5_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_5_U' read by process 'kernel_pr_kernel_pr.load_value_5_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_bipedge_U0_ap_ready & load_bipedge_U0.ap_idle & ~ap_sync_load_value_5_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_5_U0'");
                        end
                    end
                    9: begin
                        if (~load_bipedge_U0.grp_load_bipedge_Pipeline_load_bipedge_loop_fu_86.bipedge_stream_6_blk_n) begin
                            if (~bipedge_stream_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_6_U' written by process 'kernel_pr_kernel_pr.load_value_6_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_6_U' read by process 'kernel_pr_kernel_pr.load_value_6_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_bipedge_U0_ap_ready & load_bipedge_U0.ap_idle & ~ap_sync_load_value_6_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_6_U0'");
                        end
                    end
                    10: begin
                        if (~load_bipedge_U0.grp_load_bipedge_Pipeline_load_bipedge_loop_fu_86.bipedge_stream_7_blk_n) begin
                            if (~bipedge_stream_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_7_U' written by process 'kernel_pr_kernel_pr.load_value_7_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_7_U' read by process 'kernel_pr_kernel_pr.load_value_7_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_bipedge_U0_ap_ready & load_bipedge_U0.ap_idle & ~ap_sync_load_value_7_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_7_U0'");
                        end
                    end
                    0: begin
                        if (ap_sync_load_bipedge_U0_ap_ready & load_bipedge_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.entry_proc_U0'");
                        end
                    end
                    2: begin
                        if (ap_sync_load_bipedge_U0_ap_ready & load_bipedge_U0.ap_idle & ~ap_sync_load_bipedge_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge_1_U0'");
                        end
                    end
                    11: begin
                        if (ap_sync_load_bipedge_U0_ap_ready & load_bipedge_U0.ap_idle & ~ap_sync_load_value_8_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_8_U0'");
                        end
                    end
                    12: begin
                        if (ap_sync_load_bipedge_U0_ap_ready & load_bipedge_U0.ap_idle & ~ap_sync_load_value_9_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_9_U0'");
                        end
                    end
                    13: begin
                        if (ap_sync_load_bipedge_U0_ap_ready & load_bipedge_U0.ap_idle & ~ap_sync_load_value_10_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_10_U0'");
                        end
                    end
                    14: begin
                        if (ap_sync_load_bipedge_U0_ap_ready & load_bipedge_U0.ap_idle & ~ap_sync_load_value_11_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_11_U0'");
                        end
                    end
                    15: begin
                        if (ap_sync_load_bipedge_U0_ap_ready & load_bipedge_U0.ap_idle & ~ap_sync_load_value_12_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_12_U0'");
                        end
                    end
                    16: begin
                        if (ap_sync_load_bipedge_U0_ap_ready & load_bipedge_U0.ap_idle & ~ap_sync_load_value_13_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_13_U0'");
                        end
                    end
                    17: begin
                        if (ap_sync_load_bipedge_U0_ap_ready & load_bipedge_U0.ap_idle & ~ap_sync_load_value_14_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_14_U0'");
                        end
                    end
                    18: begin
                        if (ap_sync_load_bipedge_U0_ap_ready & load_bipedge_U0.ap_idle & ~ap_sync_load_value_15_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_15_U0'");
                        end
                    end
                    endcase
                end
                2 : begin
                    case(index2)
                    11: begin
                        if (~load_bipedge_1_U0.grp_load_bipedge_1_Pipeline_load_bipedge_loop_fu_86.bipedge_stream_8_blk_n) begin
                            if (~bipedge_stream_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_8_U' written by process 'kernel_pr_kernel_pr.load_value_8_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_8_U' read by process 'kernel_pr_kernel_pr.load_value_8_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_bipedge_1_U0_ap_ready & load_bipedge_1_U0.ap_idle & ~ap_sync_load_value_8_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_8_U0'");
                        end
                    end
                    12: begin
                        if (~load_bipedge_1_U0.grp_load_bipedge_1_Pipeline_load_bipedge_loop_fu_86.bipedge_stream_9_blk_n) begin
                            if (~bipedge_stream_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_9_U' written by process 'kernel_pr_kernel_pr.load_value_9_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_9_U' read by process 'kernel_pr_kernel_pr.load_value_9_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_bipedge_1_U0_ap_ready & load_bipedge_1_U0.ap_idle & ~ap_sync_load_value_9_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_9_U0'");
                        end
                    end
                    13: begin
                        if (~load_bipedge_1_U0.grp_load_bipedge_1_Pipeline_load_bipedge_loop_fu_86.bipedge_stream_10_blk_n) begin
                            if (~bipedge_stream_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_10_U' written by process 'kernel_pr_kernel_pr.load_value_10_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_10_U' read by process 'kernel_pr_kernel_pr.load_value_10_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_bipedge_1_U0_ap_ready & load_bipedge_1_U0.ap_idle & ~ap_sync_load_value_10_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_10_U0'");
                        end
                    end
                    14: begin
                        if (~load_bipedge_1_U0.grp_load_bipedge_1_Pipeline_load_bipedge_loop_fu_86.bipedge_stream_11_blk_n) begin
                            if (~bipedge_stream_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_11_U' written by process 'kernel_pr_kernel_pr.load_value_11_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_11_U' read by process 'kernel_pr_kernel_pr.load_value_11_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_bipedge_1_U0_ap_ready & load_bipedge_1_U0.ap_idle & ~ap_sync_load_value_11_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_11_U0'");
                        end
                    end
                    15: begin
                        if (~load_bipedge_1_U0.grp_load_bipedge_1_Pipeline_load_bipedge_loop_fu_86.bipedge_stream_12_blk_n) begin
                            if (~bipedge_stream_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_12_U' written by process 'kernel_pr_kernel_pr.load_value_12_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_12_U' read by process 'kernel_pr_kernel_pr.load_value_12_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_bipedge_1_U0_ap_ready & load_bipedge_1_U0.ap_idle & ~ap_sync_load_value_12_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_12_U0'");
                        end
                    end
                    16: begin
                        if (~load_bipedge_1_U0.grp_load_bipedge_1_Pipeline_load_bipedge_loop_fu_86.bipedge_stream_13_blk_n) begin
                            if (~bipedge_stream_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_13_U' written by process 'kernel_pr_kernel_pr.load_value_13_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_13_U' read by process 'kernel_pr_kernel_pr.load_value_13_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_bipedge_1_U0_ap_ready & load_bipedge_1_U0.ap_idle & ~ap_sync_load_value_13_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_13_U0'");
                        end
                    end
                    17: begin
                        if (~load_bipedge_1_U0.grp_load_bipedge_1_Pipeline_load_bipedge_loop_fu_86.bipedge_stream_14_blk_n) begin
                            if (~bipedge_stream_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_14_U' written by process 'kernel_pr_kernel_pr.load_value_14_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_14_U' read by process 'kernel_pr_kernel_pr.load_value_14_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_bipedge_1_U0_ap_ready & load_bipedge_1_U0.ap_idle & ~ap_sync_load_value_14_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_14_U0'");
                        end
                    end
                    18: begin
                        if (~load_bipedge_1_U0.grp_load_bipedge_1_Pipeline_load_bipedge_loop_fu_86.bipedge_stream_15_blk_n) begin
                            if (~bipedge_stream_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_15_U' written by process 'kernel_pr_kernel_pr.load_value_15_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_15_U' read by process 'kernel_pr_kernel_pr.load_value_15_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_bipedge_1_U0_ap_ready & load_bipedge_1_U0.ap_idle & ~ap_sync_load_value_15_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_15_U0'");
                        end
                    end
                    0: begin
                        if (ap_sync_load_bipedge_1_U0_ap_ready & load_bipedge_1_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.entry_proc_U0'");
                        end
                    end
                    1: begin
                        if (ap_sync_load_bipedge_1_U0_ap_ready & load_bipedge_1_U0.ap_idle & ~ap_sync_load_bipedge_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge_U0'");
                        end
                    end
                    3: begin
                        if (ap_sync_load_bipedge_1_U0_ap_ready & load_bipedge_1_U0.ap_idle & ~ap_sync_load_value_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_U0'");
                        end
                    end
                    4: begin
                        if (ap_sync_load_bipedge_1_U0_ap_ready & load_bipedge_1_U0.ap_idle & ~ap_sync_load_value_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_1_U0'");
                        end
                    end
                    5: begin
                        if (ap_sync_load_bipedge_1_U0_ap_ready & load_bipedge_1_U0.ap_idle & ~ap_sync_load_value_2_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_2_U0'");
                        end
                    end
                    6: begin
                        if (ap_sync_load_bipedge_1_U0_ap_ready & load_bipedge_1_U0.ap_idle & ~ap_sync_load_value_3_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_3_U0'");
                        end
                    end
                    7: begin
                        if (ap_sync_load_bipedge_1_U0_ap_ready & load_bipedge_1_U0.ap_idle & ~ap_sync_load_value_4_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_4_U0'");
                        end
                    end
                    8: begin
                        if (ap_sync_load_bipedge_1_U0_ap_ready & load_bipedge_1_U0.ap_idle & ~ap_sync_load_value_5_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_5_U0'");
                        end
                    end
                    9: begin
                        if (ap_sync_load_bipedge_1_U0_ap_ready & load_bipedge_1_U0.ap_idle & ~ap_sync_load_value_6_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_6_U0'");
                        end
                    end
                    10: begin
                        if (ap_sync_load_bipedge_1_U0_ap_ready & load_bipedge_1_U0.ap_idle & ~ap_sync_load_value_7_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_7_U0'");
                        end
                    end
                    endcase
                end
                3 : begin
                    case(index2)
                    1: begin
                        if (~load_value_U0.grp_load_value_Pipeline_load_value_fu_71.bipedge_stream_0_blk_n) begin
                            if (~bipedge_stream_0_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_0_U' written by process 'kernel_pr_kernel_pr.load_bipedge_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_0_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_0_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_0_U' read by process 'kernel_pr_kernel_pr.load_bipedge_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_0_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value_U0_ap_ready & load_value_U0.ap_idle & ~ap_sync_load_bipedge_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge_U0'");
                        end
                    end
                    19: begin
                        if (~load_value_U0.value_stream_0_blk_n) begin
                            if (~value_stream_0_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_0_U' written by process 'kernel_pr_kernel_pr.write_back_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_0_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_0_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_0_U' read by process 'kernel_pr_kernel_pr.write_back_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_0_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    0: begin
                        if (ap_sync_load_value_U0_ap_ready & load_value_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.entry_proc_U0'");
                        end
                    end
                    2: begin
                        if (ap_sync_load_value_U0_ap_ready & load_value_U0.ap_idle & ~ap_sync_load_bipedge_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge_1_U0'");
                        end
                    end
                    4: begin
                        if (ap_sync_load_value_U0_ap_ready & load_value_U0.ap_idle & ~ap_sync_load_value_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_1_U0'");
                        end
                    end
                    5: begin
                        if (ap_sync_load_value_U0_ap_ready & load_value_U0.ap_idle & ~ap_sync_load_value_2_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_2_U0'");
                        end
                    end
                    6: begin
                        if (ap_sync_load_value_U0_ap_ready & load_value_U0.ap_idle & ~ap_sync_load_value_3_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_3_U0'");
                        end
                    end
                    7: begin
                        if (ap_sync_load_value_U0_ap_ready & load_value_U0.ap_idle & ~ap_sync_load_value_4_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_4_U0'");
                        end
                    end
                    8: begin
                        if (ap_sync_load_value_U0_ap_ready & load_value_U0.ap_idle & ~ap_sync_load_value_5_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_5_U0'");
                        end
                    end
                    9: begin
                        if (ap_sync_load_value_U0_ap_ready & load_value_U0.ap_idle & ~ap_sync_load_value_6_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_6_U0'");
                        end
                    end
                    10: begin
                        if (ap_sync_load_value_U0_ap_ready & load_value_U0.ap_idle & ~ap_sync_load_value_7_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_7_U0'");
                        end
                    end
                    11: begin
                        if (ap_sync_load_value_U0_ap_ready & load_value_U0.ap_idle & ~ap_sync_load_value_8_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_8_U0'");
                        end
                    end
                    12: begin
                        if (ap_sync_load_value_U0_ap_ready & load_value_U0.ap_idle & ~ap_sync_load_value_9_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_9_U0'");
                        end
                    end
                    13: begin
                        if (ap_sync_load_value_U0_ap_ready & load_value_U0.ap_idle & ~ap_sync_load_value_10_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_10_U0'");
                        end
                    end
                    14: begin
                        if (ap_sync_load_value_U0_ap_ready & load_value_U0.ap_idle & ~ap_sync_load_value_11_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_11_U0'");
                        end
                    end
                    15: begin
                        if (ap_sync_load_value_U0_ap_ready & load_value_U0.ap_idle & ~ap_sync_load_value_12_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_12_U0'");
                        end
                    end
                    16: begin
                        if (ap_sync_load_value_U0_ap_ready & load_value_U0.ap_idle & ~ap_sync_load_value_13_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_13_U0'");
                        end
                    end
                    17: begin
                        if (ap_sync_load_value_U0_ap_ready & load_value_U0.ap_idle & ~ap_sync_load_value_14_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_14_U0'");
                        end
                    end
                    18: begin
                        if (ap_sync_load_value_U0_ap_ready & load_value_U0.ap_idle & ~ap_sync_load_value_15_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_15_U0'");
                        end
                    end
                    endcase
                end
                4 : begin
                    case(index2)
                    1: begin
                        if (~load_value_1_U0.grp_load_value_1_Pipeline_load_value_fu_71.bipedge_stream_1_blk_n) begin
                            if (~bipedge_stream_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_1_U' written by process 'kernel_pr_kernel_pr.load_bipedge_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_1_U' read by process 'kernel_pr_kernel_pr.load_bipedge_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value_1_U0_ap_ready & load_value_1_U0.ap_idle & ~ap_sync_load_bipedge_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge_U0'");
                        end
                    end
                    20: begin
                        if (~load_value_1_U0.value_stream_1_blk_n) begin
                            if (~value_stream_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_1_U' written by process 'kernel_pr_kernel_pr.write_back_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_1_U' read by process 'kernel_pr_kernel_pr.write_back_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    0: begin
                        if (ap_sync_load_value_1_U0_ap_ready & load_value_1_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.entry_proc_U0'");
                        end
                    end
                    2: begin
                        if (ap_sync_load_value_1_U0_ap_ready & load_value_1_U0.ap_idle & ~ap_sync_load_bipedge_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge_1_U0'");
                        end
                    end
                    3: begin
                        if (ap_sync_load_value_1_U0_ap_ready & load_value_1_U0.ap_idle & ~ap_sync_load_value_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_U0'");
                        end
                    end
                    5: begin
                        if (ap_sync_load_value_1_U0_ap_ready & load_value_1_U0.ap_idle & ~ap_sync_load_value_2_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_2_U0'");
                        end
                    end
                    6: begin
                        if (ap_sync_load_value_1_U0_ap_ready & load_value_1_U0.ap_idle & ~ap_sync_load_value_3_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_3_U0'");
                        end
                    end
                    7: begin
                        if (ap_sync_load_value_1_U0_ap_ready & load_value_1_U0.ap_idle & ~ap_sync_load_value_4_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_4_U0'");
                        end
                    end
                    8: begin
                        if (ap_sync_load_value_1_U0_ap_ready & load_value_1_U0.ap_idle & ~ap_sync_load_value_5_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_5_U0'");
                        end
                    end
                    9: begin
                        if (ap_sync_load_value_1_U0_ap_ready & load_value_1_U0.ap_idle & ~ap_sync_load_value_6_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_6_U0'");
                        end
                    end
                    10: begin
                        if (ap_sync_load_value_1_U0_ap_ready & load_value_1_U0.ap_idle & ~ap_sync_load_value_7_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_7_U0'");
                        end
                    end
                    11: begin
                        if (ap_sync_load_value_1_U0_ap_ready & load_value_1_U0.ap_idle & ~ap_sync_load_value_8_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_8_U0'");
                        end
                    end
                    12: begin
                        if (ap_sync_load_value_1_U0_ap_ready & load_value_1_U0.ap_idle & ~ap_sync_load_value_9_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_9_U0'");
                        end
                    end
                    13: begin
                        if (ap_sync_load_value_1_U0_ap_ready & load_value_1_U0.ap_idle & ~ap_sync_load_value_10_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_10_U0'");
                        end
                    end
                    14: begin
                        if (ap_sync_load_value_1_U0_ap_ready & load_value_1_U0.ap_idle & ~ap_sync_load_value_11_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_11_U0'");
                        end
                    end
                    15: begin
                        if (ap_sync_load_value_1_U0_ap_ready & load_value_1_U0.ap_idle & ~ap_sync_load_value_12_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_12_U0'");
                        end
                    end
                    16: begin
                        if (ap_sync_load_value_1_U0_ap_ready & load_value_1_U0.ap_idle & ~ap_sync_load_value_13_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_13_U0'");
                        end
                    end
                    17: begin
                        if (ap_sync_load_value_1_U0_ap_ready & load_value_1_U0.ap_idle & ~ap_sync_load_value_14_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_14_U0'");
                        end
                    end
                    18: begin
                        if (ap_sync_load_value_1_U0_ap_ready & load_value_1_U0.ap_idle & ~ap_sync_load_value_15_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_15_U0'");
                        end
                    end
                    endcase
                end
                5 : begin
                    case(index2)
                    1: begin
                        if (~load_value_2_U0.grp_load_value_2_Pipeline_load_value_fu_71.bipedge_stream_2_blk_n) begin
                            if (~bipedge_stream_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_2_U' written by process 'kernel_pr_kernel_pr.load_bipedge_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_2_U' read by process 'kernel_pr_kernel_pr.load_bipedge_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value_2_U0_ap_ready & load_value_2_U0.ap_idle & ~ap_sync_load_bipedge_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge_U0'");
                        end
                    end
                    21: begin
                        if (~load_value_2_U0.value_stream_2_blk_n) begin
                            if (~value_stream_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_2_U' written by process 'kernel_pr_kernel_pr.write_back_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_2_U' read by process 'kernel_pr_kernel_pr.write_back_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    0: begin
                        if (ap_sync_load_value_2_U0_ap_ready & load_value_2_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.entry_proc_U0'");
                        end
                    end
                    2: begin
                        if (ap_sync_load_value_2_U0_ap_ready & load_value_2_U0.ap_idle & ~ap_sync_load_bipedge_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge_1_U0'");
                        end
                    end
                    3: begin
                        if (ap_sync_load_value_2_U0_ap_ready & load_value_2_U0.ap_idle & ~ap_sync_load_value_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_U0'");
                        end
                    end
                    4: begin
                        if (ap_sync_load_value_2_U0_ap_ready & load_value_2_U0.ap_idle & ~ap_sync_load_value_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_1_U0'");
                        end
                    end
                    6: begin
                        if (ap_sync_load_value_2_U0_ap_ready & load_value_2_U0.ap_idle & ~ap_sync_load_value_3_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_3_U0'");
                        end
                    end
                    7: begin
                        if (ap_sync_load_value_2_U0_ap_ready & load_value_2_U0.ap_idle & ~ap_sync_load_value_4_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_4_U0'");
                        end
                    end
                    8: begin
                        if (ap_sync_load_value_2_U0_ap_ready & load_value_2_U0.ap_idle & ~ap_sync_load_value_5_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_5_U0'");
                        end
                    end
                    9: begin
                        if (ap_sync_load_value_2_U0_ap_ready & load_value_2_U0.ap_idle & ~ap_sync_load_value_6_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_6_U0'");
                        end
                    end
                    10: begin
                        if (ap_sync_load_value_2_U0_ap_ready & load_value_2_U0.ap_idle & ~ap_sync_load_value_7_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_7_U0'");
                        end
                    end
                    11: begin
                        if (ap_sync_load_value_2_U0_ap_ready & load_value_2_U0.ap_idle & ~ap_sync_load_value_8_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_8_U0'");
                        end
                    end
                    12: begin
                        if (ap_sync_load_value_2_U0_ap_ready & load_value_2_U0.ap_idle & ~ap_sync_load_value_9_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_9_U0'");
                        end
                    end
                    13: begin
                        if (ap_sync_load_value_2_U0_ap_ready & load_value_2_U0.ap_idle & ~ap_sync_load_value_10_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_10_U0'");
                        end
                    end
                    14: begin
                        if (ap_sync_load_value_2_U0_ap_ready & load_value_2_U0.ap_idle & ~ap_sync_load_value_11_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_11_U0'");
                        end
                    end
                    15: begin
                        if (ap_sync_load_value_2_U0_ap_ready & load_value_2_U0.ap_idle & ~ap_sync_load_value_12_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_12_U0'");
                        end
                    end
                    16: begin
                        if (ap_sync_load_value_2_U0_ap_ready & load_value_2_U0.ap_idle & ~ap_sync_load_value_13_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_13_U0'");
                        end
                    end
                    17: begin
                        if (ap_sync_load_value_2_U0_ap_ready & load_value_2_U0.ap_idle & ~ap_sync_load_value_14_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_14_U0'");
                        end
                    end
                    18: begin
                        if (ap_sync_load_value_2_U0_ap_ready & load_value_2_U0.ap_idle & ~ap_sync_load_value_15_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_15_U0'");
                        end
                    end
                    endcase
                end
                6 : begin
                    case(index2)
                    1: begin
                        if (~load_value_3_U0.grp_load_value_3_Pipeline_load_value_fu_71.bipedge_stream_3_blk_n) begin
                            if (~bipedge_stream_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_3_U' written by process 'kernel_pr_kernel_pr.load_bipedge_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_3_U' read by process 'kernel_pr_kernel_pr.load_bipedge_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value_3_U0_ap_ready & load_value_3_U0.ap_idle & ~ap_sync_load_bipedge_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge_U0'");
                        end
                    end
                    22: begin
                        if (~load_value_3_U0.value_stream_3_blk_n) begin
                            if (~value_stream_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_3_U' written by process 'kernel_pr_kernel_pr.write_back_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_3_U' read by process 'kernel_pr_kernel_pr.write_back_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    0: begin
                        if (ap_sync_load_value_3_U0_ap_ready & load_value_3_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.entry_proc_U0'");
                        end
                    end
                    2: begin
                        if (ap_sync_load_value_3_U0_ap_ready & load_value_3_U0.ap_idle & ~ap_sync_load_bipedge_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge_1_U0'");
                        end
                    end
                    3: begin
                        if (ap_sync_load_value_3_U0_ap_ready & load_value_3_U0.ap_idle & ~ap_sync_load_value_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_U0'");
                        end
                    end
                    4: begin
                        if (ap_sync_load_value_3_U0_ap_ready & load_value_3_U0.ap_idle & ~ap_sync_load_value_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_1_U0'");
                        end
                    end
                    5: begin
                        if (ap_sync_load_value_3_U0_ap_ready & load_value_3_U0.ap_idle & ~ap_sync_load_value_2_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_2_U0'");
                        end
                    end
                    7: begin
                        if (ap_sync_load_value_3_U0_ap_ready & load_value_3_U0.ap_idle & ~ap_sync_load_value_4_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_4_U0'");
                        end
                    end
                    8: begin
                        if (ap_sync_load_value_3_U0_ap_ready & load_value_3_U0.ap_idle & ~ap_sync_load_value_5_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_5_U0'");
                        end
                    end
                    9: begin
                        if (ap_sync_load_value_3_U0_ap_ready & load_value_3_U0.ap_idle & ~ap_sync_load_value_6_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_6_U0'");
                        end
                    end
                    10: begin
                        if (ap_sync_load_value_3_U0_ap_ready & load_value_3_U0.ap_idle & ~ap_sync_load_value_7_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_7_U0'");
                        end
                    end
                    11: begin
                        if (ap_sync_load_value_3_U0_ap_ready & load_value_3_U0.ap_idle & ~ap_sync_load_value_8_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_8_U0'");
                        end
                    end
                    12: begin
                        if (ap_sync_load_value_3_U0_ap_ready & load_value_3_U0.ap_idle & ~ap_sync_load_value_9_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_9_U0'");
                        end
                    end
                    13: begin
                        if (ap_sync_load_value_3_U0_ap_ready & load_value_3_U0.ap_idle & ~ap_sync_load_value_10_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_10_U0'");
                        end
                    end
                    14: begin
                        if (ap_sync_load_value_3_U0_ap_ready & load_value_3_U0.ap_idle & ~ap_sync_load_value_11_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_11_U0'");
                        end
                    end
                    15: begin
                        if (ap_sync_load_value_3_U0_ap_ready & load_value_3_U0.ap_idle & ~ap_sync_load_value_12_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_12_U0'");
                        end
                    end
                    16: begin
                        if (ap_sync_load_value_3_U0_ap_ready & load_value_3_U0.ap_idle & ~ap_sync_load_value_13_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_13_U0'");
                        end
                    end
                    17: begin
                        if (ap_sync_load_value_3_U0_ap_ready & load_value_3_U0.ap_idle & ~ap_sync_load_value_14_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_14_U0'");
                        end
                    end
                    18: begin
                        if (ap_sync_load_value_3_U0_ap_ready & load_value_3_U0.ap_idle & ~ap_sync_load_value_15_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_15_U0'");
                        end
                    end
                    endcase
                end
                7 : begin
                    case(index2)
                    1: begin
                        if (~load_value_4_U0.grp_load_value_4_Pipeline_load_value_fu_71.bipedge_stream_4_blk_n) begin
                            if (~bipedge_stream_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_4_U' written by process 'kernel_pr_kernel_pr.load_bipedge_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_4_U' read by process 'kernel_pr_kernel_pr.load_bipedge_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value_4_U0_ap_ready & load_value_4_U0.ap_idle & ~ap_sync_load_bipedge_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge_U0'");
                        end
                    end
                    23: begin
                        if (~load_value_4_U0.value_stream_4_blk_n) begin
                            if (~value_stream_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_4_U' written by process 'kernel_pr_kernel_pr.write_back_4_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_4_U' read by process 'kernel_pr_kernel_pr.write_back_4_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    0: begin
                        if (ap_sync_load_value_4_U0_ap_ready & load_value_4_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.entry_proc_U0'");
                        end
                    end
                    2: begin
                        if (ap_sync_load_value_4_U0_ap_ready & load_value_4_U0.ap_idle & ~ap_sync_load_bipedge_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge_1_U0'");
                        end
                    end
                    3: begin
                        if (ap_sync_load_value_4_U0_ap_ready & load_value_4_U0.ap_idle & ~ap_sync_load_value_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_U0'");
                        end
                    end
                    4: begin
                        if (ap_sync_load_value_4_U0_ap_ready & load_value_4_U0.ap_idle & ~ap_sync_load_value_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_1_U0'");
                        end
                    end
                    5: begin
                        if (ap_sync_load_value_4_U0_ap_ready & load_value_4_U0.ap_idle & ~ap_sync_load_value_2_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_2_U0'");
                        end
                    end
                    6: begin
                        if (ap_sync_load_value_4_U0_ap_ready & load_value_4_U0.ap_idle & ~ap_sync_load_value_3_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_3_U0'");
                        end
                    end
                    8: begin
                        if (ap_sync_load_value_4_U0_ap_ready & load_value_4_U0.ap_idle & ~ap_sync_load_value_5_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_5_U0'");
                        end
                    end
                    9: begin
                        if (ap_sync_load_value_4_U0_ap_ready & load_value_4_U0.ap_idle & ~ap_sync_load_value_6_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_6_U0'");
                        end
                    end
                    10: begin
                        if (ap_sync_load_value_4_U0_ap_ready & load_value_4_U0.ap_idle & ~ap_sync_load_value_7_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_7_U0'");
                        end
                    end
                    11: begin
                        if (ap_sync_load_value_4_U0_ap_ready & load_value_4_U0.ap_idle & ~ap_sync_load_value_8_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_8_U0'");
                        end
                    end
                    12: begin
                        if (ap_sync_load_value_4_U0_ap_ready & load_value_4_U0.ap_idle & ~ap_sync_load_value_9_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_9_U0'");
                        end
                    end
                    13: begin
                        if (ap_sync_load_value_4_U0_ap_ready & load_value_4_U0.ap_idle & ~ap_sync_load_value_10_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_10_U0'");
                        end
                    end
                    14: begin
                        if (ap_sync_load_value_4_U0_ap_ready & load_value_4_U0.ap_idle & ~ap_sync_load_value_11_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_11_U0'");
                        end
                    end
                    15: begin
                        if (ap_sync_load_value_4_U0_ap_ready & load_value_4_U0.ap_idle & ~ap_sync_load_value_12_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_12_U0'");
                        end
                    end
                    16: begin
                        if (ap_sync_load_value_4_U0_ap_ready & load_value_4_U0.ap_idle & ~ap_sync_load_value_13_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_13_U0'");
                        end
                    end
                    17: begin
                        if (ap_sync_load_value_4_U0_ap_ready & load_value_4_U0.ap_idle & ~ap_sync_load_value_14_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_14_U0'");
                        end
                    end
                    18: begin
                        if (ap_sync_load_value_4_U0_ap_ready & load_value_4_U0.ap_idle & ~ap_sync_load_value_15_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_15_U0'");
                        end
                    end
                    endcase
                end
                8 : begin
                    case(index2)
                    1: begin
                        if (~load_value_5_U0.grp_load_value_5_Pipeline_load_value_fu_71.bipedge_stream_5_blk_n) begin
                            if (~bipedge_stream_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_5_U' written by process 'kernel_pr_kernel_pr.load_bipedge_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_5_U' read by process 'kernel_pr_kernel_pr.load_bipedge_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value_5_U0_ap_ready & load_value_5_U0.ap_idle & ~ap_sync_load_bipedge_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge_U0'");
                        end
                    end
                    24: begin
                        if (~load_value_5_U0.value_stream_5_blk_n) begin
                            if (~value_stream_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_5_U' written by process 'kernel_pr_kernel_pr.write_back_5_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_5_U' read by process 'kernel_pr_kernel_pr.write_back_5_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    0: begin
                        if (ap_sync_load_value_5_U0_ap_ready & load_value_5_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.entry_proc_U0'");
                        end
                    end
                    2: begin
                        if (ap_sync_load_value_5_U0_ap_ready & load_value_5_U0.ap_idle & ~ap_sync_load_bipedge_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge_1_U0'");
                        end
                    end
                    3: begin
                        if (ap_sync_load_value_5_U0_ap_ready & load_value_5_U0.ap_idle & ~ap_sync_load_value_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_U0'");
                        end
                    end
                    4: begin
                        if (ap_sync_load_value_5_U0_ap_ready & load_value_5_U0.ap_idle & ~ap_sync_load_value_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_1_U0'");
                        end
                    end
                    5: begin
                        if (ap_sync_load_value_5_U0_ap_ready & load_value_5_U0.ap_idle & ~ap_sync_load_value_2_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_2_U0'");
                        end
                    end
                    6: begin
                        if (ap_sync_load_value_5_U0_ap_ready & load_value_5_U0.ap_idle & ~ap_sync_load_value_3_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_3_U0'");
                        end
                    end
                    7: begin
                        if (ap_sync_load_value_5_U0_ap_ready & load_value_5_U0.ap_idle & ~ap_sync_load_value_4_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_4_U0'");
                        end
                    end
                    9: begin
                        if (ap_sync_load_value_5_U0_ap_ready & load_value_5_U0.ap_idle & ~ap_sync_load_value_6_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_6_U0'");
                        end
                    end
                    10: begin
                        if (ap_sync_load_value_5_U0_ap_ready & load_value_5_U0.ap_idle & ~ap_sync_load_value_7_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_7_U0'");
                        end
                    end
                    11: begin
                        if (ap_sync_load_value_5_U0_ap_ready & load_value_5_U0.ap_idle & ~ap_sync_load_value_8_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_8_U0'");
                        end
                    end
                    12: begin
                        if (ap_sync_load_value_5_U0_ap_ready & load_value_5_U0.ap_idle & ~ap_sync_load_value_9_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_9_U0'");
                        end
                    end
                    13: begin
                        if (ap_sync_load_value_5_U0_ap_ready & load_value_5_U0.ap_idle & ~ap_sync_load_value_10_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_10_U0'");
                        end
                    end
                    14: begin
                        if (ap_sync_load_value_5_U0_ap_ready & load_value_5_U0.ap_idle & ~ap_sync_load_value_11_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_11_U0'");
                        end
                    end
                    15: begin
                        if (ap_sync_load_value_5_U0_ap_ready & load_value_5_U0.ap_idle & ~ap_sync_load_value_12_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_12_U0'");
                        end
                    end
                    16: begin
                        if (ap_sync_load_value_5_U0_ap_ready & load_value_5_U0.ap_idle & ~ap_sync_load_value_13_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_13_U0'");
                        end
                    end
                    17: begin
                        if (ap_sync_load_value_5_U0_ap_ready & load_value_5_U0.ap_idle & ~ap_sync_load_value_14_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_14_U0'");
                        end
                    end
                    18: begin
                        if (ap_sync_load_value_5_U0_ap_ready & load_value_5_U0.ap_idle & ~ap_sync_load_value_15_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_15_U0'");
                        end
                    end
                    endcase
                end
                9 : begin
                    case(index2)
                    1: begin
                        if (~load_value_6_U0.grp_load_value_6_Pipeline_load_value_fu_71.bipedge_stream_6_blk_n) begin
                            if (~bipedge_stream_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_6_U' written by process 'kernel_pr_kernel_pr.load_bipedge_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_6_U' read by process 'kernel_pr_kernel_pr.load_bipedge_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value_6_U0_ap_ready & load_value_6_U0.ap_idle & ~ap_sync_load_bipedge_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge_U0'");
                        end
                    end
                    25: begin
                        if (~load_value_6_U0.value_stream_6_blk_n) begin
                            if (~value_stream_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_6_U' written by process 'kernel_pr_kernel_pr.write_back_6_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_6_U' read by process 'kernel_pr_kernel_pr.write_back_6_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    0: begin
                        if (ap_sync_load_value_6_U0_ap_ready & load_value_6_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.entry_proc_U0'");
                        end
                    end
                    2: begin
                        if (ap_sync_load_value_6_U0_ap_ready & load_value_6_U0.ap_idle & ~ap_sync_load_bipedge_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge_1_U0'");
                        end
                    end
                    3: begin
                        if (ap_sync_load_value_6_U0_ap_ready & load_value_6_U0.ap_idle & ~ap_sync_load_value_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_U0'");
                        end
                    end
                    4: begin
                        if (ap_sync_load_value_6_U0_ap_ready & load_value_6_U0.ap_idle & ~ap_sync_load_value_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_1_U0'");
                        end
                    end
                    5: begin
                        if (ap_sync_load_value_6_U0_ap_ready & load_value_6_U0.ap_idle & ~ap_sync_load_value_2_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_2_U0'");
                        end
                    end
                    6: begin
                        if (ap_sync_load_value_6_U0_ap_ready & load_value_6_U0.ap_idle & ~ap_sync_load_value_3_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_3_U0'");
                        end
                    end
                    7: begin
                        if (ap_sync_load_value_6_U0_ap_ready & load_value_6_U0.ap_idle & ~ap_sync_load_value_4_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_4_U0'");
                        end
                    end
                    8: begin
                        if (ap_sync_load_value_6_U0_ap_ready & load_value_6_U0.ap_idle & ~ap_sync_load_value_5_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_5_U0'");
                        end
                    end
                    10: begin
                        if (ap_sync_load_value_6_U0_ap_ready & load_value_6_U0.ap_idle & ~ap_sync_load_value_7_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_7_U0'");
                        end
                    end
                    11: begin
                        if (ap_sync_load_value_6_U0_ap_ready & load_value_6_U0.ap_idle & ~ap_sync_load_value_8_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_8_U0'");
                        end
                    end
                    12: begin
                        if (ap_sync_load_value_6_U0_ap_ready & load_value_6_U0.ap_idle & ~ap_sync_load_value_9_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_9_U0'");
                        end
                    end
                    13: begin
                        if (ap_sync_load_value_6_U0_ap_ready & load_value_6_U0.ap_idle & ~ap_sync_load_value_10_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_10_U0'");
                        end
                    end
                    14: begin
                        if (ap_sync_load_value_6_U0_ap_ready & load_value_6_U0.ap_idle & ~ap_sync_load_value_11_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_11_U0'");
                        end
                    end
                    15: begin
                        if (ap_sync_load_value_6_U0_ap_ready & load_value_6_U0.ap_idle & ~ap_sync_load_value_12_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_12_U0'");
                        end
                    end
                    16: begin
                        if (ap_sync_load_value_6_U0_ap_ready & load_value_6_U0.ap_idle & ~ap_sync_load_value_13_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_13_U0'");
                        end
                    end
                    17: begin
                        if (ap_sync_load_value_6_U0_ap_ready & load_value_6_U0.ap_idle & ~ap_sync_load_value_14_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_14_U0'");
                        end
                    end
                    18: begin
                        if (ap_sync_load_value_6_U0_ap_ready & load_value_6_U0.ap_idle & ~ap_sync_load_value_15_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_15_U0'");
                        end
                    end
                    endcase
                end
                10 : begin
                    case(index2)
                    1: begin
                        if (~load_value_7_U0.grp_load_value_7_Pipeline_load_value_fu_71.bipedge_stream_7_blk_n) begin
                            if (~bipedge_stream_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_7_U' written by process 'kernel_pr_kernel_pr.load_bipedge_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_7_U' read by process 'kernel_pr_kernel_pr.load_bipedge_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value_7_U0_ap_ready & load_value_7_U0.ap_idle & ~ap_sync_load_bipedge_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge_U0'");
                        end
                    end
                    26: begin
                        if (~load_value_7_U0.value_stream_7_blk_n) begin
                            if (~value_stream_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_7_U' written by process 'kernel_pr_kernel_pr.write_back_7_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_7_U' read by process 'kernel_pr_kernel_pr.write_back_7_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    0: begin
                        if (ap_sync_load_value_7_U0_ap_ready & load_value_7_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.entry_proc_U0'");
                        end
                    end
                    2: begin
                        if (ap_sync_load_value_7_U0_ap_ready & load_value_7_U0.ap_idle & ~ap_sync_load_bipedge_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge_1_U0'");
                        end
                    end
                    3: begin
                        if (ap_sync_load_value_7_U0_ap_ready & load_value_7_U0.ap_idle & ~ap_sync_load_value_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_U0'");
                        end
                    end
                    4: begin
                        if (ap_sync_load_value_7_U0_ap_ready & load_value_7_U0.ap_idle & ~ap_sync_load_value_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_1_U0'");
                        end
                    end
                    5: begin
                        if (ap_sync_load_value_7_U0_ap_ready & load_value_7_U0.ap_idle & ~ap_sync_load_value_2_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_2_U0'");
                        end
                    end
                    6: begin
                        if (ap_sync_load_value_7_U0_ap_ready & load_value_7_U0.ap_idle & ~ap_sync_load_value_3_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_3_U0'");
                        end
                    end
                    7: begin
                        if (ap_sync_load_value_7_U0_ap_ready & load_value_7_U0.ap_idle & ~ap_sync_load_value_4_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_4_U0'");
                        end
                    end
                    8: begin
                        if (ap_sync_load_value_7_U0_ap_ready & load_value_7_U0.ap_idle & ~ap_sync_load_value_5_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_5_U0'");
                        end
                    end
                    9: begin
                        if (ap_sync_load_value_7_U0_ap_ready & load_value_7_U0.ap_idle & ~ap_sync_load_value_6_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_6_U0'");
                        end
                    end
                    11: begin
                        if (ap_sync_load_value_7_U0_ap_ready & load_value_7_U0.ap_idle & ~ap_sync_load_value_8_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_8_U0'");
                        end
                    end
                    12: begin
                        if (ap_sync_load_value_7_U0_ap_ready & load_value_7_U0.ap_idle & ~ap_sync_load_value_9_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_9_U0'");
                        end
                    end
                    13: begin
                        if (ap_sync_load_value_7_U0_ap_ready & load_value_7_U0.ap_idle & ~ap_sync_load_value_10_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_10_U0'");
                        end
                    end
                    14: begin
                        if (ap_sync_load_value_7_U0_ap_ready & load_value_7_U0.ap_idle & ~ap_sync_load_value_11_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_11_U0'");
                        end
                    end
                    15: begin
                        if (ap_sync_load_value_7_U0_ap_ready & load_value_7_U0.ap_idle & ~ap_sync_load_value_12_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_12_U0'");
                        end
                    end
                    16: begin
                        if (ap_sync_load_value_7_U0_ap_ready & load_value_7_U0.ap_idle & ~ap_sync_load_value_13_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_13_U0'");
                        end
                    end
                    17: begin
                        if (ap_sync_load_value_7_U0_ap_ready & load_value_7_U0.ap_idle & ~ap_sync_load_value_14_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_14_U0'");
                        end
                    end
                    18: begin
                        if (ap_sync_load_value_7_U0_ap_ready & load_value_7_U0.ap_idle & ~ap_sync_load_value_15_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_15_U0'");
                        end
                    end
                    endcase
                end
                11 : begin
                    case(index2)
                    2: begin
                        if (~load_value_8_U0.grp_load_value_8_Pipeline_load_value_fu_71.bipedge_stream_8_blk_n) begin
                            if (~bipedge_stream_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_8_U' written by process 'kernel_pr_kernel_pr.load_bipedge_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_8_U' read by process 'kernel_pr_kernel_pr.load_bipedge_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value_8_U0_ap_ready & load_value_8_U0.ap_idle & ~ap_sync_load_bipedge_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge_1_U0'");
                        end
                    end
                    27: begin
                        if (~load_value_8_U0.value_stream_8_blk_n) begin
                            if (~value_stream_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_8_U' written by process 'kernel_pr_kernel_pr.write_back_8_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_8_U' read by process 'kernel_pr_kernel_pr.write_back_8_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    0: begin
                        if (ap_sync_load_value_8_U0_ap_ready & load_value_8_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.entry_proc_U0'");
                        end
                    end
                    1: begin
                        if (ap_sync_load_value_8_U0_ap_ready & load_value_8_U0.ap_idle & ~ap_sync_load_bipedge_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge_U0'");
                        end
                    end
                    3: begin
                        if (ap_sync_load_value_8_U0_ap_ready & load_value_8_U0.ap_idle & ~ap_sync_load_value_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_U0'");
                        end
                    end
                    4: begin
                        if (ap_sync_load_value_8_U0_ap_ready & load_value_8_U0.ap_idle & ~ap_sync_load_value_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_1_U0'");
                        end
                    end
                    5: begin
                        if (ap_sync_load_value_8_U0_ap_ready & load_value_8_U0.ap_idle & ~ap_sync_load_value_2_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_2_U0'");
                        end
                    end
                    6: begin
                        if (ap_sync_load_value_8_U0_ap_ready & load_value_8_U0.ap_idle & ~ap_sync_load_value_3_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_3_U0'");
                        end
                    end
                    7: begin
                        if (ap_sync_load_value_8_U0_ap_ready & load_value_8_U0.ap_idle & ~ap_sync_load_value_4_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_4_U0'");
                        end
                    end
                    8: begin
                        if (ap_sync_load_value_8_U0_ap_ready & load_value_8_U0.ap_idle & ~ap_sync_load_value_5_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_5_U0'");
                        end
                    end
                    9: begin
                        if (ap_sync_load_value_8_U0_ap_ready & load_value_8_U0.ap_idle & ~ap_sync_load_value_6_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_6_U0'");
                        end
                    end
                    10: begin
                        if (ap_sync_load_value_8_U0_ap_ready & load_value_8_U0.ap_idle & ~ap_sync_load_value_7_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_7_U0'");
                        end
                    end
                    12: begin
                        if (ap_sync_load_value_8_U0_ap_ready & load_value_8_U0.ap_idle & ~ap_sync_load_value_9_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_9_U0'");
                        end
                    end
                    13: begin
                        if (ap_sync_load_value_8_U0_ap_ready & load_value_8_U0.ap_idle & ~ap_sync_load_value_10_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_10_U0'");
                        end
                    end
                    14: begin
                        if (ap_sync_load_value_8_U0_ap_ready & load_value_8_U0.ap_idle & ~ap_sync_load_value_11_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_11_U0'");
                        end
                    end
                    15: begin
                        if (ap_sync_load_value_8_U0_ap_ready & load_value_8_U0.ap_idle & ~ap_sync_load_value_12_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_12_U0'");
                        end
                    end
                    16: begin
                        if (ap_sync_load_value_8_U0_ap_ready & load_value_8_U0.ap_idle & ~ap_sync_load_value_13_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_13_U0'");
                        end
                    end
                    17: begin
                        if (ap_sync_load_value_8_U0_ap_ready & load_value_8_U0.ap_idle & ~ap_sync_load_value_14_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_14_U0'");
                        end
                    end
                    18: begin
                        if (ap_sync_load_value_8_U0_ap_ready & load_value_8_U0.ap_idle & ~ap_sync_load_value_15_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_15_U0'");
                        end
                    end
                    endcase
                end
                12 : begin
                    case(index2)
                    2: begin
                        if (~load_value_9_U0.grp_load_value_9_Pipeline_load_value_fu_71.bipedge_stream_9_blk_n) begin
                            if (~bipedge_stream_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_9_U' written by process 'kernel_pr_kernel_pr.load_bipedge_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_9_U' read by process 'kernel_pr_kernel_pr.load_bipedge_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value_9_U0_ap_ready & load_value_9_U0.ap_idle & ~ap_sync_load_bipedge_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge_1_U0'");
                        end
                    end
                    28: begin
                        if (~load_value_9_U0.value_stream_9_blk_n) begin
                            if (~value_stream_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_9_U' written by process 'kernel_pr_kernel_pr.write_back_9_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_9_U' read by process 'kernel_pr_kernel_pr.write_back_9_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    0: begin
                        if (ap_sync_load_value_9_U0_ap_ready & load_value_9_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.entry_proc_U0'");
                        end
                    end
                    1: begin
                        if (ap_sync_load_value_9_U0_ap_ready & load_value_9_U0.ap_idle & ~ap_sync_load_bipedge_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge_U0'");
                        end
                    end
                    3: begin
                        if (ap_sync_load_value_9_U0_ap_ready & load_value_9_U0.ap_idle & ~ap_sync_load_value_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_U0'");
                        end
                    end
                    4: begin
                        if (ap_sync_load_value_9_U0_ap_ready & load_value_9_U0.ap_idle & ~ap_sync_load_value_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_1_U0'");
                        end
                    end
                    5: begin
                        if (ap_sync_load_value_9_U0_ap_ready & load_value_9_U0.ap_idle & ~ap_sync_load_value_2_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_2_U0'");
                        end
                    end
                    6: begin
                        if (ap_sync_load_value_9_U0_ap_ready & load_value_9_U0.ap_idle & ~ap_sync_load_value_3_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_3_U0'");
                        end
                    end
                    7: begin
                        if (ap_sync_load_value_9_U0_ap_ready & load_value_9_U0.ap_idle & ~ap_sync_load_value_4_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_4_U0'");
                        end
                    end
                    8: begin
                        if (ap_sync_load_value_9_U0_ap_ready & load_value_9_U0.ap_idle & ~ap_sync_load_value_5_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_5_U0'");
                        end
                    end
                    9: begin
                        if (ap_sync_load_value_9_U0_ap_ready & load_value_9_U0.ap_idle & ~ap_sync_load_value_6_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_6_U0'");
                        end
                    end
                    10: begin
                        if (ap_sync_load_value_9_U0_ap_ready & load_value_9_U0.ap_idle & ~ap_sync_load_value_7_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_7_U0'");
                        end
                    end
                    11: begin
                        if (ap_sync_load_value_9_U0_ap_ready & load_value_9_U0.ap_idle & ~ap_sync_load_value_8_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_8_U0'");
                        end
                    end
                    13: begin
                        if (ap_sync_load_value_9_U0_ap_ready & load_value_9_U0.ap_idle & ~ap_sync_load_value_10_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_10_U0'");
                        end
                    end
                    14: begin
                        if (ap_sync_load_value_9_U0_ap_ready & load_value_9_U0.ap_idle & ~ap_sync_load_value_11_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_11_U0'");
                        end
                    end
                    15: begin
                        if (ap_sync_load_value_9_U0_ap_ready & load_value_9_U0.ap_idle & ~ap_sync_load_value_12_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_12_U0'");
                        end
                    end
                    16: begin
                        if (ap_sync_load_value_9_U0_ap_ready & load_value_9_U0.ap_idle & ~ap_sync_load_value_13_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_13_U0'");
                        end
                    end
                    17: begin
                        if (ap_sync_load_value_9_U0_ap_ready & load_value_9_U0.ap_idle & ~ap_sync_load_value_14_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_14_U0'");
                        end
                    end
                    18: begin
                        if (ap_sync_load_value_9_U0_ap_ready & load_value_9_U0.ap_idle & ~ap_sync_load_value_15_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_15_U0'");
                        end
                    end
                    endcase
                end
                13 : begin
                    case(index2)
                    2: begin
                        if (~load_value_10_U0.grp_load_value_10_Pipeline_load_value_fu_71.bipedge_stream_10_blk_n) begin
                            if (~bipedge_stream_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_10_U' written by process 'kernel_pr_kernel_pr.load_bipedge_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_10_U' read by process 'kernel_pr_kernel_pr.load_bipedge_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value_10_U0_ap_ready & load_value_10_U0.ap_idle & ~ap_sync_load_bipedge_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge_1_U0'");
                        end
                    end
                    29: begin
                        if (~load_value_10_U0.value_stream_10_blk_n) begin
                            if (~value_stream_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_10_U' written by process 'kernel_pr_kernel_pr.write_back_10_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_10_U' read by process 'kernel_pr_kernel_pr.write_back_10_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    0: begin
                        if (ap_sync_load_value_10_U0_ap_ready & load_value_10_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.entry_proc_U0'");
                        end
                    end
                    1: begin
                        if (ap_sync_load_value_10_U0_ap_ready & load_value_10_U0.ap_idle & ~ap_sync_load_bipedge_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge_U0'");
                        end
                    end
                    3: begin
                        if (ap_sync_load_value_10_U0_ap_ready & load_value_10_U0.ap_idle & ~ap_sync_load_value_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_U0'");
                        end
                    end
                    4: begin
                        if (ap_sync_load_value_10_U0_ap_ready & load_value_10_U0.ap_idle & ~ap_sync_load_value_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_1_U0'");
                        end
                    end
                    5: begin
                        if (ap_sync_load_value_10_U0_ap_ready & load_value_10_U0.ap_idle & ~ap_sync_load_value_2_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_2_U0'");
                        end
                    end
                    6: begin
                        if (ap_sync_load_value_10_U0_ap_ready & load_value_10_U0.ap_idle & ~ap_sync_load_value_3_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_3_U0'");
                        end
                    end
                    7: begin
                        if (ap_sync_load_value_10_U0_ap_ready & load_value_10_U0.ap_idle & ~ap_sync_load_value_4_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_4_U0'");
                        end
                    end
                    8: begin
                        if (ap_sync_load_value_10_U0_ap_ready & load_value_10_U0.ap_idle & ~ap_sync_load_value_5_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_5_U0'");
                        end
                    end
                    9: begin
                        if (ap_sync_load_value_10_U0_ap_ready & load_value_10_U0.ap_idle & ~ap_sync_load_value_6_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_6_U0'");
                        end
                    end
                    10: begin
                        if (ap_sync_load_value_10_U0_ap_ready & load_value_10_U0.ap_idle & ~ap_sync_load_value_7_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_7_U0'");
                        end
                    end
                    11: begin
                        if (ap_sync_load_value_10_U0_ap_ready & load_value_10_U0.ap_idle & ~ap_sync_load_value_8_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_8_U0'");
                        end
                    end
                    12: begin
                        if (ap_sync_load_value_10_U0_ap_ready & load_value_10_U0.ap_idle & ~ap_sync_load_value_9_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_9_U0'");
                        end
                    end
                    14: begin
                        if (ap_sync_load_value_10_U0_ap_ready & load_value_10_U0.ap_idle & ~ap_sync_load_value_11_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_11_U0'");
                        end
                    end
                    15: begin
                        if (ap_sync_load_value_10_U0_ap_ready & load_value_10_U0.ap_idle & ~ap_sync_load_value_12_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_12_U0'");
                        end
                    end
                    16: begin
                        if (ap_sync_load_value_10_U0_ap_ready & load_value_10_U0.ap_idle & ~ap_sync_load_value_13_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_13_U0'");
                        end
                    end
                    17: begin
                        if (ap_sync_load_value_10_U0_ap_ready & load_value_10_U0.ap_idle & ~ap_sync_load_value_14_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_14_U0'");
                        end
                    end
                    18: begin
                        if (ap_sync_load_value_10_U0_ap_ready & load_value_10_U0.ap_idle & ~ap_sync_load_value_15_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_15_U0'");
                        end
                    end
                    endcase
                end
                14 : begin
                    case(index2)
                    2: begin
                        if (~load_value_11_U0.grp_load_value_11_Pipeline_load_value_fu_71.bipedge_stream_11_blk_n) begin
                            if (~bipedge_stream_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_11_U' written by process 'kernel_pr_kernel_pr.load_bipedge_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_11_U' read by process 'kernel_pr_kernel_pr.load_bipedge_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value_11_U0_ap_ready & load_value_11_U0.ap_idle & ~ap_sync_load_bipedge_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge_1_U0'");
                        end
                    end
                    30: begin
                        if (~load_value_11_U0.value_stream_11_blk_n) begin
                            if (~value_stream_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_11_U' written by process 'kernel_pr_kernel_pr.write_back_11_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_11_U' read by process 'kernel_pr_kernel_pr.write_back_11_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    0: begin
                        if (ap_sync_load_value_11_U0_ap_ready & load_value_11_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.entry_proc_U0'");
                        end
                    end
                    1: begin
                        if (ap_sync_load_value_11_U0_ap_ready & load_value_11_U0.ap_idle & ~ap_sync_load_bipedge_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge_U0'");
                        end
                    end
                    3: begin
                        if (ap_sync_load_value_11_U0_ap_ready & load_value_11_U0.ap_idle & ~ap_sync_load_value_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_U0'");
                        end
                    end
                    4: begin
                        if (ap_sync_load_value_11_U0_ap_ready & load_value_11_U0.ap_idle & ~ap_sync_load_value_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_1_U0'");
                        end
                    end
                    5: begin
                        if (ap_sync_load_value_11_U0_ap_ready & load_value_11_U0.ap_idle & ~ap_sync_load_value_2_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_2_U0'");
                        end
                    end
                    6: begin
                        if (ap_sync_load_value_11_U0_ap_ready & load_value_11_U0.ap_idle & ~ap_sync_load_value_3_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_3_U0'");
                        end
                    end
                    7: begin
                        if (ap_sync_load_value_11_U0_ap_ready & load_value_11_U0.ap_idle & ~ap_sync_load_value_4_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_4_U0'");
                        end
                    end
                    8: begin
                        if (ap_sync_load_value_11_U0_ap_ready & load_value_11_U0.ap_idle & ~ap_sync_load_value_5_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_5_U0'");
                        end
                    end
                    9: begin
                        if (ap_sync_load_value_11_U0_ap_ready & load_value_11_U0.ap_idle & ~ap_sync_load_value_6_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_6_U0'");
                        end
                    end
                    10: begin
                        if (ap_sync_load_value_11_U0_ap_ready & load_value_11_U0.ap_idle & ~ap_sync_load_value_7_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_7_U0'");
                        end
                    end
                    11: begin
                        if (ap_sync_load_value_11_U0_ap_ready & load_value_11_U0.ap_idle & ~ap_sync_load_value_8_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_8_U0'");
                        end
                    end
                    12: begin
                        if (ap_sync_load_value_11_U0_ap_ready & load_value_11_U0.ap_idle & ~ap_sync_load_value_9_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_9_U0'");
                        end
                    end
                    13: begin
                        if (ap_sync_load_value_11_U0_ap_ready & load_value_11_U0.ap_idle & ~ap_sync_load_value_10_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_10_U0'");
                        end
                    end
                    15: begin
                        if (ap_sync_load_value_11_U0_ap_ready & load_value_11_U0.ap_idle & ~ap_sync_load_value_12_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_12_U0'");
                        end
                    end
                    16: begin
                        if (ap_sync_load_value_11_U0_ap_ready & load_value_11_U0.ap_idle & ~ap_sync_load_value_13_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_13_U0'");
                        end
                    end
                    17: begin
                        if (ap_sync_load_value_11_U0_ap_ready & load_value_11_U0.ap_idle & ~ap_sync_load_value_14_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_14_U0'");
                        end
                    end
                    18: begin
                        if (ap_sync_load_value_11_U0_ap_ready & load_value_11_U0.ap_idle & ~ap_sync_load_value_15_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_15_U0'");
                        end
                    end
                    endcase
                end
                15 : begin
                    case(index2)
                    2: begin
                        if (~load_value_12_U0.grp_load_value_12_Pipeline_load_value_fu_71.bipedge_stream_12_blk_n) begin
                            if (~bipedge_stream_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_12_U' written by process 'kernel_pr_kernel_pr.load_bipedge_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_12_U' read by process 'kernel_pr_kernel_pr.load_bipedge_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value_12_U0_ap_ready & load_value_12_U0.ap_idle & ~ap_sync_load_bipedge_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge_1_U0'");
                        end
                    end
                    31: begin
                        if (~load_value_12_U0.value_stream_12_blk_n) begin
                            if (~value_stream_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_12_U' written by process 'kernel_pr_kernel_pr.write_back_12_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_12_U' read by process 'kernel_pr_kernel_pr.write_back_12_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    0: begin
                        if (ap_sync_load_value_12_U0_ap_ready & load_value_12_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.entry_proc_U0'");
                        end
                    end
                    1: begin
                        if (ap_sync_load_value_12_U0_ap_ready & load_value_12_U0.ap_idle & ~ap_sync_load_bipedge_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge_U0'");
                        end
                    end
                    3: begin
                        if (ap_sync_load_value_12_U0_ap_ready & load_value_12_U0.ap_idle & ~ap_sync_load_value_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_U0'");
                        end
                    end
                    4: begin
                        if (ap_sync_load_value_12_U0_ap_ready & load_value_12_U0.ap_idle & ~ap_sync_load_value_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_1_U0'");
                        end
                    end
                    5: begin
                        if (ap_sync_load_value_12_U0_ap_ready & load_value_12_U0.ap_idle & ~ap_sync_load_value_2_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_2_U0'");
                        end
                    end
                    6: begin
                        if (ap_sync_load_value_12_U0_ap_ready & load_value_12_U0.ap_idle & ~ap_sync_load_value_3_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_3_U0'");
                        end
                    end
                    7: begin
                        if (ap_sync_load_value_12_U0_ap_ready & load_value_12_U0.ap_idle & ~ap_sync_load_value_4_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_4_U0'");
                        end
                    end
                    8: begin
                        if (ap_sync_load_value_12_U0_ap_ready & load_value_12_U0.ap_idle & ~ap_sync_load_value_5_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_5_U0'");
                        end
                    end
                    9: begin
                        if (ap_sync_load_value_12_U0_ap_ready & load_value_12_U0.ap_idle & ~ap_sync_load_value_6_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_6_U0'");
                        end
                    end
                    10: begin
                        if (ap_sync_load_value_12_U0_ap_ready & load_value_12_U0.ap_idle & ~ap_sync_load_value_7_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_7_U0'");
                        end
                    end
                    11: begin
                        if (ap_sync_load_value_12_U0_ap_ready & load_value_12_U0.ap_idle & ~ap_sync_load_value_8_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_8_U0'");
                        end
                    end
                    12: begin
                        if (ap_sync_load_value_12_U0_ap_ready & load_value_12_U0.ap_idle & ~ap_sync_load_value_9_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_9_U0'");
                        end
                    end
                    13: begin
                        if (ap_sync_load_value_12_U0_ap_ready & load_value_12_U0.ap_idle & ~ap_sync_load_value_10_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_10_U0'");
                        end
                    end
                    14: begin
                        if (ap_sync_load_value_12_U0_ap_ready & load_value_12_U0.ap_idle & ~ap_sync_load_value_11_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_11_U0'");
                        end
                    end
                    16: begin
                        if (ap_sync_load_value_12_U0_ap_ready & load_value_12_U0.ap_idle & ~ap_sync_load_value_13_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_13_U0'");
                        end
                    end
                    17: begin
                        if (ap_sync_load_value_12_U0_ap_ready & load_value_12_U0.ap_idle & ~ap_sync_load_value_14_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_14_U0'");
                        end
                    end
                    18: begin
                        if (ap_sync_load_value_12_U0_ap_ready & load_value_12_U0.ap_idle & ~ap_sync_load_value_15_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_15_U0'");
                        end
                    end
                    endcase
                end
                16 : begin
                    case(index2)
                    2: begin
                        if (~load_value_13_U0.grp_load_value_13_Pipeline_load_value_fu_71.bipedge_stream_13_blk_n) begin
                            if (~bipedge_stream_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_13_U' written by process 'kernel_pr_kernel_pr.load_bipedge_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_13_U' read by process 'kernel_pr_kernel_pr.load_bipedge_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value_13_U0_ap_ready & load_value_13_U0.ap_idle & ~ap_sync_load_bipedge_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge_1_U0'");
                        end
                    end
                    32: begin
                        if (~load_value_13_U0.value_stream_13_blk_n) begin
                            if (~value_stream_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_13_U' written by process 'kernel_pr_kernel_pr.write_back_13_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_13_U' read by process 'kernel_pr_kernel_pr.write_back_13_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    0: begin
                        if (ap_sync_load_value_13_U0_ap_ready & load_value_13_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.entry_proc_U0'");
                        end
                    end
                    1: begin
                        if (ap_sync_load_value_13_U0_ap_ready & load_value_13_U0.ap_idle & ~ap_sync_load_bipedge_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge_U0'");
                        end
                    end
                    3: begin
                        if (ap_sync_load_value_13_U0_ap_ready & load_value_13_U0.ap_idle & ~ap_sync_load_value_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_U0'");
                        end
                    end
                    4: begin
                        if (ap_sync_load_value_13_U0_ap_ready & load_value_13_U0.ap_idle & ~ap_sync_load_value_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_1_U0'");
                        end
                    end
                    5: begin
                        if (ap_sync_load_value_13_U0_ap_ready & load_value_13_U0.ap_idle & ~ap_sync_load_value_2_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_2_U0'");
                        end
                    end
                    6: begin
                        if (ap_sync_load_value_13_U0_ap_ready & load_value_13_U0.ap_idle & ~ap_sync_load_value_3_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_3_U0'");
                        end
                    end
                    7: begin
                        if (ap_sync_load_value_13_U0_ap_ready & load_value_13_U0.ap_idle & ~ap_sync_load_value_4_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_4_U0'");
                        end
                    end
                    8: begin
                        if (ap_sync_load_value_13_U0_ap_ready & load_value_13_U0.ap_idle & ~ap_sync_load_value_5_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_5_U0'");
                        end
                    end
                    9: begin
                        if (ap_sync_load_value_13_U0_ap_ready & load_value_13_U0.ap_idle & ~ap_sync_load_value_6_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_6_U0'");
                        end
                    end
                    10: begin
                        if (ap_sync_load_value_13_U0_ap_ready & load_value_13_U0.ap_idle & ~ap_sync_load_value_7_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_7_U0'");
                        end
                    end
                    11: begin
                        if (ap_sync_load_value_13_U0_ap_ready & load_value_13_U0.ap_idle & ~ap_sync_load_value_8_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_8_U0'");
                        end
                    end
                    12: begin
                        if (ap_sync_load_value_13_U0_ap_ready & load_value_13_U0.ap_idle & ~ap_sync_load_value_9_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_9_U0'");
                        end
                    end
                    13: begin
                        if (ap_sync_load_value_13_U0_ap_ready & load_value_13_U0.ap_idle & ~ap_sync_load_value_10_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_10_U0'");
                        end
                    end
                    14: begin
                        if (ap_sync_load_value_13_U0_ap_ready & load_value_13_U0.ap_idle & ~ap_sync_load_value_11_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_11_U0'");
                        end
                    end
                    15: begin
                        if (ap_sync_load_value_13_U0_ap_ready & load_value_13_U0.ap_idle & ~ap_sync_load_value_12_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_12_U0'");
                        end
                    end
                    17: begin
                        if (ap_sync_load_value_13_U0_ap_ready & load_value_13_U0.ap_idle & ~ap_sync_load_value_14_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_14_U0'");
                        end
                    end
                    18: begin
                        if (ap_sync_load_value_13_U0_ap_ready & load_value_13_U0.ap_idle & ~ap_sync_load_value_15_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_15_U0'");
                        end
                    end
                    endcase
                end
                17 : begin
                    case(index2)
                    2: begin
                        if (~load_value_14_U0.grp_load_value_14_Pipeline_load_value_fu_71.bipedge_stream_14_blk_n) begin
                            if (~bipedge_stream_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_14_U' written by process 'kernel_pr_kernel_pr.load_bipedge_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_14_U' read by process 'kernel_pr_kernel_pr.load_bipedge_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value_14_U0_ap_ready & load_value_14_U0.ap_idle & ~ap_sync_load_bipedge_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge_1_U0'");
                        end
                    end
                    33: begin
                        if (~load_value_14_U0.value_stream_14_blk_n) begin
                            if (~value_stream_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_14_U' written by process 'kernel_pr_kernel_pr.write_back_14_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_14_U' read by process 'kernel_pr_kernel_pr.write_back_14_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    0: begin
                        if (ap_sync_load_value_14_U0_ap_ready & load_value_14_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.entry_proc_U0'");
                        end
                    end
                    1: begin
                        if (ap_sync_load_value_14_U0_ap_ready & load_value_14_U0.ap_idle & ~ap_sync_load_bipedge_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge_U0'");
                        end
                    end
                    3: begin
                        if (ap_sync_load_value_14_U0_ap_ready & load_value_14_U0.ap_idle & ~ap_sync_load_value_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_U0'");
                        end
                    end
                    4: begin
                        if (ap_sync_load_value_14_U0_ap_ready & load_value_14_U0.ap_idle & ~ap_sync_load_value_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_1_U0'");
                        end
                    end
                    5: begin
                        if (ap_sync_load_value_14_U0_ap_ready & load_value_14_U0.ap_idle & ~ap_sync_load_value_2_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_2_U0'");
                        end
                    end
                    6: begin
                        if (ap_sync_load_value_14_U0_ap_ready & load_value_14_U0.ap_idle & ~ap_sync_load_value_3_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_3_U0'");
                        end
                    end
                    7: begin
                        if (ap_sync_load_value_14_U0_ap_ready & load_value_14_U0.ap_idle & ~ap_sync_load_value_4_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_4_U0'");
                        end
                    end
                    8: begin
                        if (ap_sync_load_value_14_U0_ap_ready & load_value_14_U0.ap_idle & ~ap_sync_load_value_5_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_5_U0'");
                        end
                    end
                    9: begin
                        if (ap_sync_load_value_14_U0_ap_ready & load_value_14_U0.ap_idle & ~ap_sync_load_value_6_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_6_U0'");
                        end
                    end
                    10: begin
                        if (ap_sync_load_value_14_U0_ap_ready & load_value_14_U0.ap_idle & ~ap_sync_load_value_7_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_7_U0'");
                        end
                    end
                    11: begin
                        if (ap_sync_load_value_14_U0_ap_ready & load_value_14_U0.ap_idle & ~ap_sync_load_value_8_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_8_U0'");
                        end
                    end
                    12: begin
                        if (ap_sync_load_value_14_U0_ap_ready & load_value_14_U0.ap_idle & ~ap_sync_load_value_9_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_9_U0'");
                        end
                    end
                    13: begin
                        if (ap_sync_load_value_14_U0_ap_ready & load_value_14_U0.ap_idle & ~ap_sync_load_value_10_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_10_U0'");
                        end
                    end
                    14: begin
                        if (ap_sync_load_value_14_U0_ap_ready & load_value_14_U0.ap_idle & ~ap_sync_load_value_11_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_11_U0'");
                        end
                    end
                    15: begin
                        if (ap_sync_load_value_14_U0_ap_ready & load_value_14_U0.ap_idle & ~ap_sync_load_value_12_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_12_U0'");
                        end
                    end
                    16: begin
                        if (ap_sync_load_value_14_U0_ap_ready & load_value_14_U0.ap_idle & ~ap_sync_load_value_13_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_13_U0'");
                        end
                    end
                    18: begin
                        if (ap_sync_load_value_14_U0_ap_ready & load_value_14_U0.ap_idle & ~ap_sync_load_value_15_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_15_U0'");
                        end
                    end
                    endcase
                end
                18 : begin
                    case(index2)
                    2: begin
                        if (~load_value_15_U0.grp_load_value_15_Pipeline_load_value_fu_71.bipedge_stream_15_blk_n) begin
                            if (~bipedge_stream_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_15_U' written by process 'kernel_pr_kernel_pr.load_bipedge_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_15_U' read by process 'kernel_pr_kernel_pr.load_bipedge_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value_15_U0_ap_ready & load_value_15_U0.ap_idle & ~ap_sync_load_bipedge_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge_1_U0'");
                        end
                    end
                    34: begin
                        if (~load_value_15_U0.value_stream_15_blk_n) begin
                            if (~value_stream_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_15_U' written by process 'kernel_pr_kernel_pr.write_back_15_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_15_U' read by process 'kernel_pr_kernel_pr.write_back_15_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    0: begin
                        if (ap_sync_load_value_15_U0_ap_ready & load_value_15_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.entry_proc_U0'");
                        end
                    end
                    1: begin
                        if (ap_sync_load_value_15_U0_ap_ready & load_value_15_U0.ap_idle & ~ap_sync_load_bipedge_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge_U0'");
                        end
                    end
                    3: begin
                        if (ap_sync_load_value_15_U0_ap_ready & load_value_15_U0.ap_idle & ~ap_sync_load_value_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_U0'");
                        end
                    end
                    4: begin
                        if (ap_sync_load_value_15_U0_ap_ready & load_value_15_U0.ap_idle & ~ap_sync_load_value_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_1_U0'");
                        end
                    end
                    5: begin
                        if (ap_sync_load_value_15_U0_ap_ready & load_value_15_U0.ap_idle & ~ap_sync_load_value_2_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_2_U0'");
                        end
                    end
                    6: begin
                        if (ap_sync_load_value_15_U0_ap_ready & load_value_15_U0.ap_idle & ~ap_sync_load_value_3_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_3_U0'");
                        end
                    end
                    7: begin
                        if (ap_sync_load_value_15_U0_ap_ready & load_value_15_U0.ap_idle & ~ap_sync_load_value_4_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_4_U0'");
                        end
                    end
                    8: begin
                        if (ap_sync_load_value_15_U0_ap_ready & load_value_15_U0.ap_idle & ~ap_sync_load_value_5_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_5_U0'");
                        end
                    end
                    9: begin
                        if (ap_sync_load_value_15_U0_ap_ready & load_value_15_U0.ap_idle & ~ap_sync_load_value_6_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_6_U0'");
                        end
                    end
                    10: begin
                        if (ap_sync_load_value_15_U0_ap_ready & load_value_15_U0.ap_idle & ~ap_sync_load_value_7_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_7_U0'");
                        end
                    end
                    11: begin
                        if (ap_sync_load_value_15_U0_ap_ready & load_value_15_U0.ap_idle & ~ap_sync_load_value_8_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_8_U0'");
                        end
                    end
                    12: begin
                        if (ap_sync_load_value_15_U0_ap_ready & load_value_15_U0.ap_idle & ~ap_sync_load_value_9_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_9_U0'");
                        end
                    end
                    13: begin
                        if (ap_sync_load_value_15_U0_ap_ready & load_value_15_U0.ap_idle & ~ap_sync_load_value_10_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_10_U0'");
                        end
                    end
                    14: begin
                        if (ap_sync_load_value_15_U0_ap_ready & load_value_15_U0.ap_idle & ~ap_sync_load_value_11_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_11_U0'");
                        end
                    end
                    15: begin
                        if (ap_sync_load_value_15_U0_ap_ready & load_value_15_U0.ap_idle & ~ap_sync_load_value_12_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_12_U0'");
                        end
                    end
                    16: begin
                        if (ap_sync_load_value_15_U0_ap_ready & load_value_15_U0.ap_idle & ~ap_sync_load_value_13_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_13_U0'");
                        end
                    end
                    17: begin
                        if (ap_sync_load_value_15_U0_ap_ready & load_value_15_U0.ap_idle & ~ap_sync_load_value_14_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value_14_U0'");
                        end
                    end
                    endcase
                end
                19 : begin
                    case(index2)
                    0: begin
                        if (~write_back_U0.H_blk_n) begin
                            if (~H_write0_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write0_c_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write0_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write0_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write0_c_U' read by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write0_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~write_back_U0.hyperedge_size_blk_n) begin
                            if (~hyperedge_size_c85_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c85_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c85_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c85_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c85_U' read by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c85_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back_U0_U.if_empty_n & write_back_U0.ap_idle & ~start_for_write_back_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back_U0_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0',");
                        end
                    end
                    3: begin
                        if (~write_back_U0.grp_write_back_Pipeline_write_back_loop_fu_81.value_stream_0_blk_n) begin
                            if (~value_stream_0_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_0_U' written by process 'kernel_pr_kernel_pr.load_value_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_0_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_0_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_0_U' read by process 'kernel_pr_kernel_pr.load_value_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_0_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    20: begin
                        if (ap_done_reg_0 & write_back_U0.ap_done & ~write_back_1_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_1_U0'");
                        end
                    end
                    21: begin
                        if (ap_done_reg_0 & write_back_U0.ap_done & ~write_back_2_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_2_U0'");
                        end
                    end
                    22: begin
                        if (ap_done_reg_0 & write_back_U0.ap_done & ~write_back_3_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_3_U0'");
                        end
                    end
                    23: begin
                        if (ap_done_reg_0 & write_back_U0.ap_done & ~write_back_4_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_4_U0'");
                        end
                    end
                    24: begin
                        if (ap_done_reg_0 & write_back_U0.ap_done & ~write_back_5_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_5_U0'");
                        end
                    end
                    25: begin
                        if (ap_done_reg_0 & write_back_U0.ap_done & ~write_back_6_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_6_U0'");
                        end
                    end
                    26: begin
                        if (ap_done_reg_0 & write_back_U0.ap_done & ~write_back_7_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_7_U0'");
                        end
                    end
                    27: begin
                        if (ap_done_reg_0 & write_back_U0.ap_done & ~write_back_8_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_8_U0'");
                        end
                    end
                    28: begin
                        if (ap_done_reg_0 & write_back_U0.ap_done & ~write_back_9_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_9_U0'");
                        end
                    end
                    29: begin
                        if (ap_done_reg_0 & write_back_U0.ap_done & ~write_back_10_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_10_U0'");
                        end
                    end
                    30: begin
                        if (ap_done_reg_0 & write_back_U0.ap_done & ~write_back_11_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_11_U0'");
                        end
                    end
                    31: begin
                        if (ap_done_reg_0 & write_back_U0.ap_done & ~write_back_12_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_12_U0'");
                        end
                    end
                    32: begin
                        if (ap_done_reg_0 & write_back_U0.ap_done & ~write_back_13_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_13_U0'");
                        end
                    end
                    33: begin
                        if (ap_done_reg_0 & write_back_U0.ap_done & ~write_back_14_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_14_U0'");
                        end
                    end
                    34: begin
                        if (ap_done_reg_0 & write_back_U0.ap_done & ~write_back_15_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_15_U0'");
                        end
                    end
                    endcase
                end
                20 : begin
                    case(index2)
                    0: begin
                        if (~write_back_1_U0.H_blk_n) begin
                            if (~H_write1_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write1_c_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write1_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write1_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write1_c_U' read by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write1_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~write_back_1_U0.hyperedge_size_blk_n) begin
                            if (~hyperedge_size_c84_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c84_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c84_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c84_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c84_U' read by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c84_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back_1_U0_U.if_empty_n & write_back_1_U0.ap_idle & ~start_for_write_back_1_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back_1_U0_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0',");
                        end
                    end
                    4: begin
                        if (~write_back_1_U0.grp_write_back_1_Pipeline_write_back_loop_fu_87.value_stream_1_blk_n) begin
                            if (~value_stream_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_1_U' written by process 'kernel_pr_kernel_pr.load_value_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_1_U' read by process 'kernel_pr_kernel_pr.load_value_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin
                        if (ap_done_reg_1 & write_back_1_U0.ap_done & ~write_back_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_U0'");
                        end
                    end
                    21: begin
                        if (ap_done_reg_1 & write_back_1_U0.ap_done & ~write_back_2_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_2_U0'");
                        end
                    end
                    22: begin
                        if (ap_done_reg_1 & write_back_1_U0.ap_done & ~write_back_3_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_3_U0'");
                        end
                    end
                    23: begin
                        if (ap_done_reg_1 & write_back_1_U0.ap_done & ~write_back_4_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_4_U0'");
                        end
                    end
                    24: begin
                        if (ap_done_reg_1 & write_back_1_U0.ap_done & ~write_back_5_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_5_U0'");
                        end
                    end
                    25: begin
                        if (ap_done_reg_1 & write_back_1_U0.ap_done & ~write_back_6_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_6_U0'");
                        end
                    end
                    26: begin
                        if (ap_done_reg_1 & write_back_1_U0.ap_done & ~write_back_7_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_7_U0'");
                        end
                    end
                    27: begin
                        if (ap_done_reg_1 & write_back_1_U0.ap_done & ~write_back_8_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_8_U0'");
                        end
                    end
                    28: begin
                        if (ap_done_reg_1 & write_back_1_U0.ap_done & ~write_back_9_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_9_U0'");
                        end
                    end
                    29: begin
                        if (ap_done_reg_1 & write_back_1_U0.ap_done & ~write_back_10_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_10_U0'");
                        end
                    end
                    30: begin
                        if (ap_done_reg_1 & write_back_1_U0.ap_done & ~write_back_11_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_11_U0'");
                        end
                    end
                    31: begin
                        if (ap_done_reg_1 & write_back_1_U0.ap_done & ~write_back_12_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_12_U0'");
                        end
                    end
                    32: begin
                        if (ap_done_reg_1 & write_back_1_U0.ap_done & ~write_back_13_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_13_U0'");
                        end
                    end
                    33: begin
                        if (ap_done_reg_1 & write_back_1_U0.ap_done & ~write_back_14_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_14_U0'");
                        end
                    end
                    34: begin
                        if (ap_done_reg_1 & write_back_1_U0.ap_done & ~write_back_15_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_15_U0'");
                        end
                    end
                    endcase
                end
                21 : begin
                    case(index2)
                    0: begin
                        if (~write_back_2_U0.H_blk_n) begin
                            if (~H_write2_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write2_c_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write2_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write2_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write2_c_U' read by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write2_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~write_back_2_U0.hyperedge_size_blk_n) begin
                            if (~hyperedge_size_c83_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c83_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c83_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c83_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c83_U' read by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c83_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back_2_U0_U.if_empty_n & write_back_2_U0.ap_idle & ~start_for_write_back_2_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back_2_U0_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0',");
                        end
                    end
                    5: begin
                        if (~write_back_2_U0.grp_write_back_2_Pipeline_write_back_loop_fu_81.value_stream_2_blk_n) begin
                            if (~value_stream_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_2_U' written by process 'kernel_pr_kernel_pr.load_value_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_2_U' read by process 'kernel_pr_kernel_pr.load_value_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin
                        if (ap_done_reg_2 & write_back_2_U0.ap_done & ~write_back_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_U0'");
                        end
                    end
                    20: begin
                        if (ap_done_reg_2 & write_back_2_U0.ap_done & ~write_back_1_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_1_U0'");
                        end
                    end
                    22: begin
                        if (ap_done_reg_2 & write_back_2_U0.ap_done & ~write_back_3_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_3_U0'");
                        end
                    end
                    23: begin
                        if (ap_done_reg_2 & write_back_2_U0.ap_done & ~write_back_4_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_4_U0'");
                        end
                    end
                    24: begin
                        if (ap_done_reg_2 & write_back_2_U0.ap_done & ~write_back_5_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_5_U0'");
                        end
                    end
                    25: begin
                        if (ap_done_reg_2 & write_back_2_U0.ap_done & ~write_back_6_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_6_U0'");
                        end
                    end
                    26: begin
                        if (ap_done_reg_2 & write_back_2_U0.ap_done & ~write_back_7_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_7_U0'");
                        end
                    end
                    27: begin
                        if (ap_done_reg_2 & write_back_2_U0.ap_done & ~write_back_8_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_8_U0'");
                        end
                    end
                    28: begin
                        if (ap_done_reg_2 & write_back_2_U0.ap_done & ~write_back_9_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_9_U0'");
                        end
                    end
                    29: begin
                        if (ap_done_reg_2 & write_back_2_U0.ap_done & ~write_back_10_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_10_U0'");
                        end
                    end
                    30: begin
                        if (ap_done_reg_2 & write_back_2_U0.ap_done & ~write_back_11_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_11_U0'");
                        end
                    end
                    31: begin
                        if (ap_done_reg_2 & write_back_2_U0.ap_done & ~write_back_12_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_12_U0'");
                        end
                    end
                    32: begin
                        if (ap_done_reg_2 & write_back_2_U0.ap_done & ~write_back_13_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_13_U0'");
                        end
                    end
                    33: begin
                        if (ap_done_reg_2 & write_back_2_U0.ap_done & ~write_back_14_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_14_U0'");
                        end
                    end
                    34: begin
                        if (ap_done_reg_2 & write_back_2_U0.ap_done & ~write_back_15_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_15_U0'");
                        end
                    end
                    endcase
                end
                22 : begin
                    case(index2)
                    0: begin
                        if (~write_back_3_U0.H_blk_n) begin
                            if (~H_write3_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write3_c_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write3_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write3_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write3_c_U' read by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write3_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~write_back_3_U0.hyperedge_size_blk_n) begin
                            if (~hyperedge_size_c82_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c82_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c82_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c82_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c82_U' read by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c82_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back_3_U0_U.if_empty_n & write_back_3_U0.ap_idle & ~start_for_write_back_3_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back_3_U0_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0',");
                        end
                    end
                    6: begin
                        if (~write_back_3_U0.grp_write_back_3_Pipeline_write_back_loop_fu_85.value_stream_3_blk_n) begin
                            if (~value_stream_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_3_U' written by process 'kernel_pr_kernel_pr.load_value_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_3_U' read by process 'kernel_pr_kernel_pr.load_value_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin
                        if (ap_done_reg_3 & write_back_3_U0.ap_done & ~write_back_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_U0'");
                        end
                    end
                    20: begin
                        if (ap_done_reg_3 & write_back_3_U0.ap_done & ~write_back_1_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_1_U0'");
                        end
                    end
                    21: begin
                        if (ap_done_reg_3 & write_back_3_U0.ap_done & ~write_back_2_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_2_U0'");
                        end
                    end
                    23: begin
                        if (ap_done_reg_3 & write_back_3_U0.ap_done & ~write_back_4_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_4_U0'");
                        end
                    end
                    24: begin
                        if (ap_done_reg_3 & write_back_3_U0.ap_done & ~write_back_5_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_5_U0'");
                        end
                    end
                    25: begin
                        if (ap_done_reg_3 & write_back_3_U0.ap_done & ~write_back_6_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_6_U0'");
                        end
                    end
                    26: begin
                        if (ap_done_reg_3 & write_back_3_U0.ap_done & ~write_back_7_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_7_U0'");
                        end
                    end
                    27: begin
                        if (ap_done_reg_3 & write_back_3_U0.ap_done & ~write_back_8_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_8_U0'");
                        end
                    end
                    28: begin
                        if (ap_done_reg_3 & write_back_3_U0.ap_done & ~write_back_9_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_9_U0'");
                        end
                    end
                    29: begin
                        if (ap_done_reg_3 & write_back_3_U0.ap_done & ~write_back_10_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_10_U0'");
                        end
                    end
                    30: begin
                        if (ap_done_reg_3 & write_back_3_U0.ap_done & ~write_back_11_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_11_U0'");
                        end
                    end
                    31: begin
                        if (ap_done_reg_3 & write_back_3_U0.ap_done & ~write_back_12_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_12_U0'");
                        end
                    end
                    32: begin
                        if (ap_done_reg_3 & write_back_3_U0.ap_done & ~write_back_13_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_13_U0'");
                        end
                    end
                    33: begin
                        if (ap_done_reg_3 & write_back_3_U0.ap_done & ~write_back_14_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_14_U0'");
                        end
                    end
                    34: begin
                        if (ap_done_reg_3 & write_back_3_U0.ap_done & ~write_back_15_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_15_U0'");
                        end
                    end
                    endcase
                end
                23 : begin
                    case(index2)
                    0: begin
                        if (~write_back_4_U0.H_blk_n) begin
                            if (~H_write4_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write4_c_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write4_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write4_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write4_c_U' read by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write4_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~write_back_4_U0.hyperedge_size_blk_n) begin
                            if (~hyperedge_size_c81_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c81_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c81_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c81_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c81_U' read by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c81_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back_4_U0_U.if_empty_n & write_back_4_U0.ap_idle & ~start_for_write_back_4_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back_4_U0_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0',");
                        end
                    end
                    7: begin
                        if (~write_back_4_U0.grp_write_back_4_Pipeline_write_back_loop_fu_81.value_stream_4_blk_n) begin
                            if (~value_stream_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_4_U' written by process 'kernel_pr_kernel_pr.load_value_4_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_4_U' read by process 'kernel_pr_kernel_pr.load_value_4_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin
                        if (ap_done_reg_4 & write_back_4_U0.ap_done & ~write_back_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_U0'");
                        end
                    end
                    20: begin
                        if (ap_done_reg_4 & write_back_4_U0.ap_done & ~write_back_1_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_1_U0'");
                        end
                    end
                    21: begin
                        if (ap_done_reg_4 & write_back_4_U0.ap_done & ~write_back_2_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_2_U0'");
                        end
                    end
                    22: begin
                        if (ap_done_reg_4 & write_back_4_U0.ap_done & ~write_back_3_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_3_U0'");
                        end
                    end
                    24: begin
                        if (ap_done_reg_4 & write_back_4_U0.ap_done & ~write_back_5_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_5_U0'");
                        end
                    end
                    25: begin
                        if (ap_done_reg_4 & write_back_4_U0.ap_done & ~write_back_6_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_6_U0'");
                        end
                    end
                    26: begin
                        if (ap_done_reg_4 & write_back_4_U0.ap_done & ~write_back_7_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_7_U0'");
                        end
                    end
                    27: begin
                        if (ap_done_reg_4 & write_back_4_U0.ap_done & ~write_back_8_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_8_U0'");
                        end
                    end
                    28: begin
                        if (ap_done_reg_4 & write_back_4_U0.ap_done & ~write_back_9_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_9_U0'");
                        end
                    end
                    29: begin
                        if (ap_done_reg_4 & write_back_4_U0.ap_done & ~write_back_10_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_10_U0'");
                        end
                    end
                    30: begin
                        if (ap_done_reg_4 & write_back_4_U0.ap_done & ~write_back_11_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_11_U0'");
                        end
                    end
                    31: begin
                        if (ap_done_reg_4 & write_back_4_U0.ap_done & ~write_back_12_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_12_U0'");
                        end
                    end
                    32: begin
                        if (ap_done_reg_4 & write_back_4_U0.ap_done & ~write_back_13_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_13_U0'");
                        end
                    end
                    33: begin
                        if (ap_done_reg_4 & write_back_4_U0.ap_done & ~write_back_14_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_14_U0'");
                        end
                    end
                    34: begin
                        if (ap_done_reg_4 & write_back_4_U0.ap_done & ~write_back_15_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_15_U0'");
                        end
                    end
                    endcase
                end
                24 : begin
                    case(index2)
                    0: begin
                        if (~write_back_5_U0.H_blk_n) begin
                            if (~H_write5_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write5_c_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write5_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write5_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write5_c_U' read by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write5_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~write_back_5_U0.hyperedge_size_blk_n) begin
                            if (~hyperedge_size_c80_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c80_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c80_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c80_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c80_U' read by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c80_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back_5_U0_U.if_empty_n & write_back_5_U0.ap_idle & ~start_for_write_back_5_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back_5_U0_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0',");
                        end
                    end
                    8: begin
                        if (~write_back_5_U0.grp_write_back_5_Pipeline_write_back_loop_fu_81.value_stream_5_blk_n) begin
                            if (~value_stream_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_5_U' written by process 'kernel_pr_kernel_pr.load_value_5_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_5_U' read by process 'kernel_pr_kernel_pr.load_value_5_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin
                        if (ap_done_reg_5 & write_back_5_U0.ap_done & ~write_back_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_U0'");
                        end
                    end
                    20: begin
                        if (ap_done_reg_5 & write_back_5_U0.ap_done & ~write_back_1_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_1_U0'");
                        end
                    end
                    21: begin
                        if (ap_done_reg_5 & write_back_5_U0.ap_done & ~write_back_2_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_2_U0'");
                        end
                    end
                    22: begin
                        if (ap_done_reg_5 & write_back_5_U0.ap_done & ~write_back_3_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_3_U0'");
                        end
                    end
                    23: begin
                        if (ap_done_reg_5 & write_back_5_U0.ap_done & ~write_back_4_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_4_U0'");
                        end
                    end
                    25: begin
                        if (ap_done_reg_5 & write_back_5_U0.ap_done & ~write_back_6_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_6_U0'");
                        end
                    end
                    26: begin
                        if (ap_done_reg_5 & write_back_5_U0.ap_done & ~write_back_7_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_7_U0'");
                        end
                    end
                    27: begin
                        if (ap_done_reg_5 & write_back_5_U0.ap_done & ~write_back_8_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_8_U0'");
                        end
                    end
                    28: begin
                        if (ap_done_reg_5 & write_back_5_U0.ap_done & ~write_back_9_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_9_U0'");
                        end
                    end
                    29: begin
                        if (ap_done_reg_5 & write_back_5_U0.ap_done & ~write_back_10_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_10_U0'");
                        end
                    end
                    30: begin
                        if (ap_done_reg_5 & write_back_5_U0.ap_done & ~write_back_11_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_11_U0'");
                        end
                    end
                    31: begin
                        if (ap_done_reg_5 & write_back_5_U0.ap_done & ~write_back_12_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_12_U0'");
                        end
                    end
                    32: begin
                        if (ap_done_reg_5 & write_back_5_U0.ap_done & ~write_back_13_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_13_U0'");
                        end
                    end
                    33: begin
                        if (ap_done_reg_5 & write_back_5_U0.ap_done & ~write_back_14_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_14_U0'");
                        end
                    end
                    34: begin
                        if (ap_done_reg_5 & write_back_5_U0.ap_done & ~write_back_15_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_15_U0'");
                        end
                    end
                    endcase
                end
                25 : begin
                    case(index2)
                    0: begin
                        if (~write_back_6_U0.H_blk_n) begin
                            if (~H_write6_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write6_c_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write6_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write6_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write6_c_U' read by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write6_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~write_back_6_U0.hyperedge_size_blk_n) begin
                            if (~hyperedge_size_c79_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c79_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c79_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c79_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c79_U' read by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c79_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back_6_U0_U.if_empty_n & write_back_6_U0.ap_idle & ~start_for_write_back_6_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back_6_U0_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0',");
                        end
                    end
                    9: begin
                        if (~write_back_6_U0.grp_write_back_6_Pipeline_write_back_loop_fu_81.value_stream_6_blk_n) begin
                            if (~value_stream_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_6_U' written by process 'kernel_pr_kernel_pr.load_value_6_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_6_U' read by process 'kernel_pr_kernel_pr.load_value_6_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin
                        if (ap_done_reg_6 & write_back_6_U0.ap_done & ~write_back_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_U0'");
                        end
                    end
                    20: begin
                        if (ap_done_reg_6 & write_back_6_U0.ap_done & ~write_back_1_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_1_U0'");
                        end
                    end
                    21: begin
                        if (ap_done_reg_6 & write_back_6_U0.ap_done & ~write_back_2_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_2_U0'");
                        end
                    end
                    22: begin
                        if (ap_done_reg_6 & write_back_6_U0.ap_done & ~write_back_3_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_3_U0'");
                        end
                    end
                    23: begin
                        if (ap_done_reg_6 & write_back_6_U0.ap_done & ~write_back_4_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_4_U0'");
                        end
                    end
                    24: begin
                        if (ap_done_reg_6 & write_back_6_U0.ap_done & ~write_back_5_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_5_U0'");
                        end
                    end
                    26: begin
                        if (ap_done_reg_6 & write_back_6_U0.ap_done & ~write_back_7_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_7_U0'");
                        end
                    end
                    27: begin
                        if (ap_done_reg_6 & write_back_6_U0.ap_done & ~write_back_8_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_8_U0'");
                        end
                    end
                    28: begin
                        if (ap_done_reg_6 & write_back_6_U0.ap_done & ~write_back_9_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_9_U0'");
                        end
                    end
                    29: begin
                        if (ap_done_reg_6 & write_back_6_U0.ap_done & ~write_back_10_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_10_U0'");
                        end
                    end
                    30: begin
                        if (ap_done_reg_6 & write_back_6_U0.ap_done & ~write_back_11_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_11_U0'");
                        end
                    end
                    31: begin
                        if (ap_done_reg_6 & write_back_6_U0.ap_done & ~write_back_12_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_12_U0'");
                        end
                    end
                    32: begin
                        if (ap_done_reg_6 & write_back_6_U0.ap_done & ~write_back_13_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_13_U0'");
                        end
                    end
                    33: begin
                        if (ap_done_reg_6 & write_back_6_U0.ap_done & ~write_back_14_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_14_U0'");
                        end
                    end
                    34: begin
                        if (ap_done_reg_6 & write_back_6_U0.ap_done & ~write_back_15_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_15_U0'");
                        end
                    end
                    endcase
                end
                26 : begin
                    case(index2)
                    0: begin
                        if (~write_back_7_U0.H_blk_n) begin
                            if (~H_write7_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write7_c_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write7_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write7_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write7_c_U' read by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write7_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~write_back_7_U0.hyperedge_size_blk_n) begin
                            if (~hyperedge_size_c78_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c78_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c78_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c78_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c78_U' read by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c78_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back_7_U0_U.if_empty_n & write_back_7_U0.ap_idle & ~start_for_write_back_7_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back_7_U0_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0',");
                        end
                    end
                    10: begin
                        if (~write_back_7_U0.grp_write_back_7_Pipeline_write_back_loop_fu_83.value_stream_7_blk_n) begin
                            if (~value_stream_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_7_U' written by process 'kernel_pr_kernel_pr.load_value_7_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_7_U' read by process 'kernel_pr_kernel_pr.load_value_7_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin
                        if (ap_done_reg_7 & write_back_7_U0.ap_done & ~write_back_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_U0'");
                        end
                    end
                    20: begin
                        if (ap_done_reg_7 & write_back_7_U0.ap_done & ~write_back_1_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_1_U0'");
                        end
                    end
                    21: begin
                        if (ap_done_reg_7 & write_back_7_U0.ap_done & ~write_back_2_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_2_U0'");
                        end
                    end
                    22: begin
                        if (ap_done_reg_7 & write_back_7_U0.ap_done & ~write_back_3_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_3_U0'");
                        end
                    end
                    23: begin
                        if (ap_done_reg_7 & write_back_7_U0.ap_done & ~write_back_4_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_4_U0'");
                        end
                    end
                    24: begin
                        if (ap_done_reg_7 & write_back_7_U0.ap_done & ~write_back_5_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_5_U0'");
                        end
                    end
                    25: begin
                        if (ap_done_reg_7 & write_back_7_U0.ap_done & ~write_back_6_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_6_U0'");
                        end
                    end
                    27: begin
                        if (ap_done_reg_7 & write_back_7_U0.ap_done & ~write_back_8_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_8_U0'");
                        end
                    end
                    28: begin
                        if (ap_done_reg_7 & write_back_7_U0.ap_done & ~write_back_9_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_9_U0'");
                        end
                    end
                    29: begin
                        if (ap_done_reg_7 & write_back_7_U0.ap_done & ~write_back_10_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_10_U0'");
                        end
                    end
                    30: begin
                        if (ap_done_reg_7 & write_back_7_U0.ap_done & ~write_back_11_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_11_U0'");
                        end
                    end
                    31: begin
                        if (ap_done_reg_7 & write_back_7_U0.ap_done & ~write_back_12_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_12_U0'");
                        end
                    end
                    32: begin
                        if (ap_done_reg_7 & write_back_7_U0.ap_done & ~write_back_13_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_13_U0'");
                        end
                    end
                    33: begin
                        if (ap_done_reg_7 & write_back_7_U0.ap_done & ~write_back_14_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_14_U0'");
                        end
                    end
                    34: begin
                        if (ap_done_reg_7 & write_back_7_U0.ap_done & ~write_back_15_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_15_U0'");
                        end
                    end
                    endcase
                end
                27 : begin
                    case(index2)
                    0: begin
                        if (~write_back_8_U0.H_blk_n) begin
                            if (~H_write8_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write8_c_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write8_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write8_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write8_c_U' read by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write8_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~write_back_8_U0.hyperedge_size_blk_n) begin
                            if (~hyperedge_size_c77_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c77_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c77_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c77_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c77_U' read by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c77_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back_8_U0_U.if_empty_n & write_back_8_U0.ap_idle & ~start_for_write_back_8_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back_8_U0_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0',");
                        end
                    end
                    11: begin
                        if (~write_back_8_U0.grp_write_back_8_Pipeline_write_back_loop_fu_81.value_stream_8_blk_n) begin
                            if (~value_stream_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_8_U' written by process 'kernel_pr_kernel_pr.load_value_8_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_8_U' read by process 'kernel_pr_kernel_pr.load_value_8_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin
                        if (ap_done_reg_8 & write_back_8_U0.ap_done & ~write_back_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_U0'");
                        end
                    end
                    20: begin
                        if (ap_done_reg_8 & write_back_8_U0.ap_done & ~write_back_1_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_1_U0'");
                        end
                    end
                    21: begin
                        if (ap_done_reg_8 & write_back_8_U0.ap_done & ~write_back_2_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_2_U0'");
                        end
                    end
                    22: begin
                        if (ap_done_reg_8 & write_back_8_U0.ap_done & ~write_back_3_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_3_U0'");
                        end
                    end
                    23: begin
                        if (ap_done_reg_8 & write_back_8_U0.ap_done & ~write_back_4_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_4_U0'");
                        end
                    end
                    24: begin
                        if (ap_done_reg_8 & write_back_8_U0.ap_done & ~write_back_5_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_5_U0'");
                        end
                    end
                    25: begin
                        if (ap_done_reg_8 & write_back_8_U0.ap_done & ~write_back_6_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_6_U0'");
                        end
                    end
                    26: begin
                        if (ap_done_reg_8 & write_back_8_U0.ap_done & ~write_back_7_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_7_U0'");
                        end
                    end
                    28: begin
                        if (ap_done_reg_8 & write_back_8_U0.ap_done & ~write_back_9_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_9_U0'");
                        end
                    end
                    29: begin
                        if (ap_done_reg_8 & write_back_8_U0.ap_done & ~write_back_10_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_10_U0'");
                        end
                    end
                    30: begin
                        if (ap_done_reg_8 & write_back_8_U0.ap_done & ~write_back_11_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_11_U0'");
                        end
                    end
                    31: begin
                        if (ap_done_reg_8 & write_back_8_U0.ap_done & ~write_back_12_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_12_U0'");
                        end
                    end
                    32: begin
                        if (ap_done_reg_8 & write_back_8_U0.ap_done & ~write_back_13_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_13_U0'");
                        end
                    end
                    33: begin
                        if (ap_done_reg_8 & write_back_8_U0.ap_done & ~write_back_14_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_14_U0'");
                        end
                    end
                    34: begin
                        if (ap_done_reg_8 & write_back_8_U0.ap_done & ~write_back_15_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_15_U0'");
                        end
                    end
                    endcase
                end
                28 : begin
                    case(index2)
                    0: begin
                        if (~write_back_9_U0.H_blk_n) begin
                            if (~H_write9_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write9_c_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write9_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write9_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write9_c_U' read by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write9_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~write_back_9_U0.hyperedge_size_blk_n) begin
                            if (~hyperedge_size_c76_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c76_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c76_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c76_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c76_U' read by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c76_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back_9_U0_U.if_empty_n & write_back_9_U0.ap_idle & ~start_for_write_back_9_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back_9_U0_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0',");
                        end
                    end
                    12: begin
                        if (~write_back_9_U0.grp_write_back_9_Pipeline_write_back_loop_fu_81.value_stream_9_blk_n) begin
                            if (~value_stream_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_9_U' written by process 'kernel_pr_kernel_pr.load_value_9_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_9_U' read by process 'kernel_pr_kernel_pr.load_value_9_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin
                        if (ap_done_reg_9 & write_back_9_U0.ap_done & ~write_back_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_U0'");
                        end
                    end
                    20: begin
                        if (ap_done_reg_9 & write_back_9_U0.ap_done & ~write_back_1_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_1_U0'");
                        end
                    end
                    21: begin
                        if (ap_done_reg_9 & write_back_9_U0.ap_done & ~write_back_2_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_2_U0'");
                        end
                    end
                    22: begin
                        if (ap_done_reg_9 & write_back_9_U0.ap_done & ~write_back_3_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_3_U0'");
                        end
                    end
                    23: begin
                        if (ap_done_reg_9 & write_back_9_U0.ap_done & ~write_back_4_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_4_U0'");
                        end
                    end
                    24: begin
                        if (ap_done_reg_9 & write_back_9_U0.ap_done & ~write_back_5_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_5_U0'");
                        end
                    end
                    25: begin
                        if (ap_done_reg_9 & write_back_9_U0.ap_done & ~write_back_6_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_6_U0'");
                        end
                    end
                    26: begin
                        if (ap_done_reg_9 & write_back_9_U0.ap_done & ~write_back_7_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_7_U0'");
                        end
                    end
                    27: begin
                        if (ap_done_reg_9 & write_back_9_U0.ap_done & ~write_back_8_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_8_U0'");
                        end
                    end
                    29: begin
                        if (ap_done_reg_9 & write_back_9_U0.ap_done & ~write_back_10_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_10_U0'");
                        end
                    end
                    30: begin
                        if (ap_done_reg_9 & write_back_9_U0.ap_done & ~write_back_11_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_11_U0'");
                        end
                    end
                    31: begin
                        if (ap_done_reg_9 & write_back_9_U0.ap_done & ~write_back_12_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_12_U0'");
                        end
                    end
                    32: begin
                        if (ap_done_reg_9 & write_back_9_U0.ap_done & ~write_back_13_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_13_U0'");
                        end
                    end
                    33: begin
                        if (ap_done_reg_9 & write_back_9_U0.ap_done & ~write_back_14_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_14_U0'");
                        end
                    end
                    34: begin
                        if (ap_done_reg_9 & write_back_9_U0.ap_done & ~write_back_15_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_15_U0'");
                        end
                    end
                    endcase
                end
                29 : begin
                    case(index2)
                    0: begin
                        if (~write_back_10_U0.H_blk_n) begin
                            if (~H_write10_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write10_c_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write10_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write10_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write10_c_U' read by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write10_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~write_back_10_U0.hyperedge_size_blk_n) begin
                            if (~hyperedge_size_c75_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c75_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c75_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c75_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c75_U' read by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c75_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back_10_U0_U.if_empty_n & write_back_10_U0.ap_idle & ~start_for_write_back_10_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back_10_U0_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0',");
                        end
                    end
                    13: begin
                        if (~write_back_10_U0.grp_write_back_10_Pipeline_write_back_loop_fu_81.value_stream_10_blk_n) begin
                            if (~value_stream_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_10_U' written by process 'kernel_pr_kernel_pr.load_value_10_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_10_U' read by process 'kernel_pr_kernel_pr.load_value_10_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin
                        if (ap_done_reg_10 & write_back_10_U0.ap_done & ~write_back_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_U0'");
                        end
                    end
                    20: begin
                        if (ap_done_reg_10 & write_back_10_U0.ap_done & ~write_back_1_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_1_U0'");
                        end
                    end
                    21: begin
                        if (ap_done_reg_10 & write_back_10_U0.ap_done & ~write_back_2_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_2_U0'");
                        end
                    end
                    22: begin
                        if (ap_done_reg_10 & write_back_10_U0.ap_done & ~write_back_3_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_3_U0'");
                        end
                    end
                    23: begin
                        if (ap_done_reg_10 & write_back_10_U0.ap_done & ~write_back_4_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_4_U0'");
                        end
                    end
                    24: begin
                        if (ap_done_reg_10 & write_back_10_U0.ap_done & ~write_back_5_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_5_U0'");
                        end
                    end
                    25: begin
                        if (ap_done_reg_10 & write_back_10_U0.ap_done & ~write_back_6_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_6_U0'");
                        end
                    end
                    26: begin
                        if (ap_done_reg_10 & write_back_10_U0.ap_done & ~write_back_7_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_7_U0'");
                        end
                    end
                    27: begin
                        if (ap_done_reg_10 & write_back_10_U0.ap_done & ~write_back_8_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_8_U0'");
                        end
                    end
                    28: begin
                        if (ap_done_reg_10 & write_back_10_U0.ap_done & ~write_back_9_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_9_U0'");
                        end
                    end
                    30: begin
                        if (ap_done_reg_10 & write_back_10_U0.ap_done & ~write_back_11_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_11_U0'");
                        end
                    end
                    31: begin
                        if (ap_done_reg_10 & write_back_10_U0.ap_done & ~write_back_12_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_12_U0'");
                        end
                    end
                    32: begin
                        if (ap_done_reg_10 & write_back_10_U0.ap_done & ~write_back_13_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_13_U0'");
                        end
                    end
                    33: begin
                        if (ap_done_reg_10 & write_back_10_U0.ap_done & ~write_back_14_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_14_U0'");
                        end
                    end
                    34: begin
                        if (ap_done_reg_10 & write_back_10_U0.ap_done & ~write_back_15_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_15_U0'");
                        end
                    end
                    endcase
                end
                30 : begin
                    case(index2)
                    0: begin
                        if (~write_back_11_U0.H_blk_n) begin
                            if (~H_write11_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write11_c_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write11_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write11_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write11_c_U' read by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write11_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~write_back_11_U0.hyperedge_size_blk_n) begin
                            if (~hyperedge_size_c74_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c74_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c74_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c74_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c74_U' read by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c74_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back_11_U0_U.if_empty_n & write_back_11_U0.ap_idle & ~start_for_write_back_11_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back_11_U0_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0',");
                        end
                    end
                    14: begin
                        if (~write_back_11_U0.grp_write_back_11_Pipeline_write_back_loop_fu_81.value_stream_11_blk_n) begin
                            if (~value_stream_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_11_U' written by process 'kernel_pr_kernel_pr.load_value_11_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_11_U' read by process 'kernel_pr_kernel_pr.load_value_11_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin
                        if (ap_done_reg_11 & write_back_11_U0.ap_done & ~write_back_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_U0'");
                        end
                    end
                    20: begin
                        if (ap_done_reg_11 & write_back_11_U0.ap_done & ~write_back_1_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_1_U0'");
                        end
                    end
                    21: begin
                        if (ap_done_reg_11 & write_back_11_U0.ap_done & ~write_back_2_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_2_U0'");
                        end
                    end
                    22: begin
                        if (ap_done_reg_11 & write_back_11_U0.ap_done & ~write_back_3_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_3_U0'");
                        end
                    end
                    23: begin
                        if (ap_done_reg_11 & write_back_11_U0.ap_done & ~write_back_4_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_4_U0'");
                        end
                    end
                    24: begin
                        if (ap_done_reg_11 & write_back_11_U0.ap_done & ~write_back_5_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_5_U0'");
                        end
                    end
                    25: begin
                        if (ap_done_reg_11 & write_back_11_U0.ap_done & ~write_back_6_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_6_U0'");
                        end
                    end
                    26: begin
                        if (ap_done_reg_11 & write_back_11_U0.ap_done & ~write_back_7_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_7_U0'");
                        end
                    end
                    27: begin
                        if (ap_done_reg_11 & write_back_11_U0.ap_done & ~write_back_8_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_8_U0'");
                        end
                    end
                    28: begin
                        if (ap_done_reg_11 & write_back_11_U0.ap_done & ~write_back_9_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_9_U0'");
                        end
                    end
                    29: begin
                        if (ap_done_reg_11 & write_back_11_U0.ap_done & ~write_back_10_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_10_U0'");
                        end
                    end
                    31: begin
                        if (ap_done_reg_11 & write_back_11_U0.ap_done & ~write_back_12_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_12_U0'");
                        end
                    end
                    32: begin
                        if (ap_done_reg_11 & write_back_11_U0.ap_done & ~write_back_13_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_13_U0'");
                        end
                    end
                    33: begin
                        if (ap_done_reg_11 & write_back_11_U0.ap_done & ~write_back_14_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_14_U0'");
                        end
                    end
                    34: begin
                        if (ap_done_reg_11 & write_back_11_U0.ap_done & ~write_back_15_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_15_U0'");
                        end
                    end
                    endcase
                end
                31 : begin
                    case(index2)
                    0: begin
                        if (~write_back_12_U0.H_blk_n) begin
                            if (~H_write12_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write12_c_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write12_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write12_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write12_c_U' read by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write12_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~write_back_12_U0.hyperedge_size_blk_n) begin
                            if (~hyperedge_size_c73_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c73_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c73_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c73_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c73_U' read by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c73_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back_12_U0_U.if_empty_n & write_back_12_U0.ap_idle & ~start_for_write_back_12_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back_12_U0_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0',");
                        end
                    end
                    15: begin
                        if (~write_back_12_U0.grp_write_back_12_Pipeline_write_back_loop_fu_81.value_stream_12_blk_n) begin
                            if (~value_stream_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_12_U' written by process 'kernel_pr_kernel_pr.load_value_12_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_12_U' read by process 'kernel_pr_kernel_pr.load_value_12_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin
                        if (ap_done_reg_12 & write_back_12_U0.ap_done & ~write_back_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_U0'");
                        end
                    end
                    20: begin
                        if (ap_done_reg_12 & write_back_12_U0.ap_done & ~write_back_1_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_1_U0'");
                        end
                    end
                    21: begin
                        if (ap_done_reg_12 & write_back_12_U0.ap_done & ~write_back_2_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_2_U0'");
                        end
                    end
                    22: begin
                        if (ap_done_reg_12 & write_back_12_U0.ap_done & ~write_back_3_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_3_U0'");
                        end
                    end
                    23: begin
                        if (ap_done_reg_12 & write_back_12_U0.ap_done & ~write_back_4_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_4_U0'");
                        end
                    end
                    24: begin
                        if (ap_done_reg_12 & write_back_12_U0.ap_done & ~write_back_5_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_5_U0'");
                        end
                    end
                    25: begin
                        if (ap_done_reg_12 & write_back_12_U0.ap_done & ~write_back_6_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_6_U0'");
                        end
                    end
                    26: begin
                        if (ap_done_reg_12 & write_back_12_U0.ap_done & ~write_back_7_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_7_U0'");
                        end
                    end
                    27: begin
                        if (ap_done_reg_12 & write_back_12_U0.ap_done & ~write_back_8_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_8_U0'");
                        end
                    end
                    28: begin
                        if (ap_done_reg_12 & write_back_12_U0.ap_done & ~write_back_9_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_9_U0'");
                        end
                    end
                    29: begin
                        if (ap_done_reg_12 & write_back_12_U0.ap_done & ~write_back_10_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_10_U0'");
                        end
                    end
                    30: begin
                        if (ap_done_reg_12 & write_back_12_U0.ap_done & ~write_back_11_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_11_U0'");
                        end
                    end
                    32: begin
                        if (ap_done_reg_12 & write_back_12_U0.ap_done & ~write_back_13_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_13_U0'");
                        end
                    end
                    33: begin
                        if (ap_done_reg_12 & write_back_12_U0.ap_done & ~write_back_14_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_14_U0'");
                        end
                    end
                    34: begin
                        if (ap_done_reg_12 & write_back_12_U0.ap_done & ~write_back_15_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_15_U0'");
                        end
                    end
                    endcase
                end
                32 : begin
                    case(index2)
                    0: begin
                        if (~write_back_13_U0.H_blk_n) begin
                            if (~H_write13_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write13_c_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write13_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write13_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write13_c_U' read by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write13_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~write_back_13_U0.hyperedge_size_blk_n) begin
                            if (~hyperedge_size_c72_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c72_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c72_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c72_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c72_U' read by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c72_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back_13_U0_U.if_empty_n & write_back_13_U0.ap_idle & ~start_for_write_back_13_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back_13_U0_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0',");
                        end
                    end
                    16: begin
                        if (~write_back_13_U0.grp_write_back_13_Pipeline_write_back_loop_fu_81.value_stream_13_blk_n) begin
                            if (~value_stream_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_13_U' written by process 'kernel_pr_kernel_pr.load_value_13_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_13_U' read by process 'kernel_pr_kernel_pr.load_value_13_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin
                        if (ap_done_reg_13 & write_back_13_U0.ap_done & ~write_back_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_U0'");
                        end
                    end
                    20: begin
                        if (ap_done_reg_13 & write_back_13_U0.ap_done & ~write_back_1_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_1_U0'");
                        end
                    end
                    21: begin
                        if (ap_done_reg_13 & write_back_13_U0.ap_done & ~write_back_2_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_2_U0'");
                        end
                    end
                    22: begin
                        if (ap_done_reg_13 & write_back_13_U0.ap_done & ~write_back_3_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_3_U0'");
                        end
                    end
                    23: begin
                        if (ap_done_reg_13 & write_back_13_U0.ap_done & ~write_back_4_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_4_U0'");
                        end
                    end
                    24: begin
                        if (ap_done_reg_13 & write_back_13_U0.ap_done & ~write_back_5_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_5_U0'");
                        end
                    end
                    25: begin
                        if (ap_done_reg_13 & write_back_13_U0.ap_done & ~write_back_6_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_6_U0'");
                        end
                    end
                    26: begin
                        if (ap_done_reg_13 & write_back_13_U0.ap_done & ~write_back_7_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_7_U0'");
                        end
                    end
                    27: begin
                        if (ap_done_reg_13 & write_back_13_U0.ap_done & ~write_back_8_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_8_U0'");
                        end
                    end
                    28: begin
                        if (ap_done_reg_13 & write_back_13_U0.ap_done & ~write_back_9_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_9_U0'");
                        end
                    end
                    29: begin
                        if (ap_done_reg_13 & write_back_13_U0.ap_done & ~write_back_10_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_10_U0'");
                        end
                    end
                    30: begin
                        if (ap_done_reg_13 & write_back_13_U0.ap_done & ~write_back_11_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_11_U0'");
                        end
                    end
                    31: begin
                        if (ap_done_reg_13 & write_back_13_U0.ap_done & ~write_back_12_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_12_U0'");
                        end
                    end
                    33: begin
                        if (ap_done_reg_13 & write_back_13_U0.ap_done & ~write_back_14_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_14_U0'");
                        end
                    end
                    34: begin
                        if (ap_done_reg_13 & write_back_13_U0.ap_done & ~write_back_15_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_15_U0'");
                        end
                    end
                    endcase
                end
                33 : begin
                    case(index2)
                    0: begin
                        if (~write_back_14_U0.H_blk_n) begin
                            if (~H_write14_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write14_c_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write14_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write14_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write14_c_U' read by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write14_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~write_back_14_U0.hyperedge_size_blk_n) begin
                            if (~hyperedge_size_c71_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c71_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c71_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c71_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c71_U' read by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c71_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back_14_U0_U.if_empty_n & write_back_14_U0.ap_idle & ~start_for_write_back_14_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back_14_U0_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0',");
                        end
                    end
                    17: begin
                        if (~write_back_14_U0.grp_write_back_14_Pipeline_write_back_loop_fu_81.value_stream_14_blk_n) begin
                            if (~value_stream_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_14_U' written by process 'kernel_pr_kernel_pr.load_value_14_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_14_U' read by process 'kernel_pr_kernel_pr.load_value_14_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin
                        if (ap_done_reg_14 & write_back_14_U0.ap_done & ~write_back_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_U0'");
                        end
                    end
                    20: begin
                        if (ap_done_reg_14 & write_back_14_U0.ap_done & ~write_back_1_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_1_U0'");
                        end
                    end
                    21: begin
                        if (ap_done_reg_14 & write_back_14_U0.ap_done & ~write_back_2_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_2_U0'");
                        end
                    end
                    22: begin
                        if (ap_done_reg_14 & write_back_14_U0.ap_done & ~write_back_3_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_3_U0'");
                        end
                    end
                    23: begin
                        if (ap_done_reg_14 & write_back_14_U0.ap_done & ~write_back_4_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_4_U0'");
                        end
                    end
                    24: begin
                        if (ap_done_reg_14 & write_back_14_U0.ap_done & ~write_back_5_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_5_U0'");
                        end
                    end
                    25: begin
                        if (ap_done_reg_14 & write_back_14_U0.ap_done & ~write_back_6_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_6_U0'");
                        end
                    end
                    26: begin
                        if (ap_done_reg_14 & write_back_14_U0.ap_done & ~write_back_7_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_7_U0'");
                        end
                    end
                    27: begin
                        if (ap_done_reg_14 & write_back_14_U0.ap_done & ~write_back_8_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_8_U0'");
                        end
                    end
                    28: begin
                        if (ap_done_reg_14 & write_back_14_U0.ap_done & ~write_back_9_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_9_U0'");
                        end
                    end
                    29: begin
                        if (ap_done_reg_14 & write_back_14_U0.ap_done & ~write_back_10_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_10_U0'");
                        end
                    end
                    30: begin
                        if (ap_done_reg_14 & write_back_14_U0.ap_done & ~write_back_11_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_11_U0'");
                        end
                    end
                    31: begin
                        if (ap_done_reg_14 & write_back_14_U0.ap_done & ~write_back_12_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_12_U0'");
                        end
                    end
                    32: begin
                        if (ap_done_reg_14 & write_back_14_U0.ap_done & ~write_back_13_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_13_U0'");
                        end
                    end
                    34: begin
                        if (ap_done_reg_14 & write_back_14_U0.ap_done & ~write_back_15_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_15_U0'");
                        end
                    end
                    endcase
                end
                34 : begin
                    case(index2)
                    0: begin
                        if (~write_back_15_U0.H_blk_n) begin
                            if (~H_write15_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write15_c_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write15_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write15_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write15_c_U' read by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write15_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~write_back_15_U0.hyperedge_size_blk_n) begin
                            if (~hyperedge_size_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c_U' read by process 'kernel_pr_kernel_pr.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back_15_U0_U.if_empty_n & write_back_15_U0.ap_idle & ~start_for_write_back_15_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back_15_U0_U' written by process 'kernel_pr_kernel_pr.entry_proc_U0',");
                        end
                    end
                    18: begin
                        if (~write_back_15_U0.grp_write_back_15_Pipeline_write_back_loop_fu_77.value_stream_15_blk_n) begin
                            if (~value_stream_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_15_U' written by process 'kernel_pr_kernel_pr.load_value_15_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_15_U' read by process 'kernel_pr_kernel_pr.load_value_15_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin
                        if (ap_done_reg_15 & write_back_15_U0.ap_done & ~write_back_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_U0'");
                        end
                    end
                    20: begin
                        if (ap_done_reg_15 & write_back_15_U0.ap_done & ~write_back_1_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_1_U0'");
                        end
                    end
                    21: begin
                        if (ap_done_reg_15 & write_back_15_U0.ap_done & ~write_back_2_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_2_U0'");
                        end
                    end
                    22: begin
                        if (ap_done_reg_15 & write_back_15_U0.ap_done & ~write_back_3_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_3_U0'");
                        end
                    end
                    23: begin
                        if (ap_done_reg_15 & write_back_15_U0.ap_done & ~write_back_4_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_4_U0'");
                        end
                    end
                    24: begin
                        if (ap_done_reg_15 & write_back_15_U0.ap_done & ~write_back_5_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_5_U0'");
                        end
                    end
                    25: begin
                        if (ap_done_reg_15 & write_back_15_U0.ap_done & ~write_back_6_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_6_U0'");
                        end
                    end
                    26: begin
                        if (ap_done_reg_15 & write_back_15_U0.ap_done & ~write_back_7_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_7_U0'");
                        end
                    end
                    27: begin
                        if (ap_done_reg_15 & write_back_15_U0.ap_done & ~write_back_8_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_8_U0'");
                        end
                    end
                    28: begin
                        if (ap_done_reg_15 & write_back_15_U0.ap_done & ~write_back_9_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_9_U0'");
                        end
                    end
                    29: begin
                        if (ap_done_reg_15 & write_back_15_U0.ap_done & ~write_back_10_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_10_U0'");
                        end
                    end
                    30: begin
                        if (ap_done_reg_15 & write_back_15_U0.ap_done & ~write_back_11_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_11_U0'");
                        end
                    end
                    31: begin
                        if (ap_done_reg_15 & write_back_15_U0.ap_done & ~write_back_12_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_12_U0'");
                        end
                    end
                    32: begin
                        if (ap_done_reg_15 & write_back_15_U0.ap_done & ~write_back_13_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_13_U0'");
                        end
                    end
                    33: begin
                        if (ap_done_reg_15 & write_back_15_U0.ap_done & ~write_back_14_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back_14_U0'");
                        end
                    end
                    endcase
                end
            endcase
        end
    endtask

    // report
    initial begin : report_deadlock
        integer cycle_id;
        integer cycle_comp_id;
        integer record_time;
        wait (dl_reset == 1);
        cycle_id = 1;
        record_time = 0;
        while (1) begin
            @ (negedge dl_clock);
            case (CS_fsm)
                ST_DL_DETECTED: begin
                    cycle_comp_id = 2;
                    if (dl_detect_reg != dl_done_reg) begin
                        if (dl_done_reg == 'b0) begin
                            print_dl_head;
                            record_time = $time;
                        end
                        print_cycle_start(proc_path(origin), cycle_id);
                        cycle_id = cycle_id + 1;
                    end
                    else begin
                        print_dl_end((cycle_id - 1),record_time);
                        @(negedge dl_clock);
                        @(negedge dl_clock);
                        $finish;
                    end
                end
                ST_DL_REPORT: begin
                    if ((|(dl_in_vec)) & ~(|(dl_in_vec & origin_reg))) begin
                        print_cycle_chan_comp(dl_in_vec_reg, dl_in_vec);
                        print_cycle_proc_comp(proc_path(dl_in_vec), cycle_comp_id);
                        cycle_comp_id = cycle_comp_id + 1;
                    end
                    else begin
                        print_cycle_chan_comp(dl_in_vec_reg, dl_in_vec);
                    end
                end
            endcase
        end
    end
 
